// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition"

// DATE "08/15/2020 00:42:35"

// 
// Device: Altera 10CL025YU256C8G Package UFBGA256
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module kyogenrv_fpga (
	clk_clk,
	kyogenrv_0_counter_readdata,
	pio_0_external_connection_export,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
input 	clk_clk;
output 	[31:0] kyogenrv_0_counter_readdata;
output 	[31:0] pio_0_external_connection_export;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \pio_0|data_out[16]~q ;
wire \pio_0|data_out[17]~q ;
wire \pio_0|data_out[18]~q ;
wire \pio_0|data_out[19]~q ;
wire \pio_0|data_out[20]~q ;
wire \pio_0|data_out[21]~q ;
wire \pio_0|data_out[22]~q ;
wire \pio_0|data_out[23]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ;
wire \kyogenrv_0|krv|id_npc[0]~q ;
wire \kyogenrv_0|krv|id_npc[1]~q ;
wire \kyogenrv_0|krv|id_pc[2]~q ;
wire \kyogenrv_0|krv|id_pc[3]~q ;
wire \kyogenrv_0|krv|id_pc[4]~q ;
wire \kyogenrv_0|krv|id_pc[5]~q ;
wire \kyogenrv_0|krv|id_pc[6]~q ;
wire \kyogenrv_0|krv|id_pc[7]~q ;
wire \kyogenrv_0|krv|id_pc[8]~q ;
wire \kyogenrv_0|krv|id_pc[9]~q ;
wire \kyogenrv_0|krv|id_pc[10]~q ;
wire \kyogenrv_0|krv|id_pc[11]~q ;
wire \kyogenrv_0|krv|id_pc[12]~q ;
wire \kyogenrv_0|krv|id_pc[13]~q ;
wire \kyogenrv_0|krv|id_pc[14]~q ;
wire \kyogenrv_0|krv|id_pc[15]~q ;
wire \kyogenrv_0|krv|id_pc[16]~q ;
wire \kyogenrv_0|krv|id_pc[17]~q ;
wire \kyogenrv_0|krv|id_pc[18]~q ;
wire \kyogenrv_0|krv|id_pc[19]~q ;
wire \kyogenrv_0|krv|id_pc[20]~q ;
wire \kyogenrv_0|krv|id_pc[21]~q ;
wire \kyogenrv_0|krv|id_pc[22]~q ;
wire \kyogenrv_0|krv|id_pc[23]~q ;
wire \kyogenrv_0|krv|id_pc[24]~q ;
wire \kyogenrv_0|krv|id_pc[25]~q ;
wire \kyogenrv_0|krv|id_pc[26]~q ;
wire \kyogenrv_0|krv|id_pc[27]~q ;
wire \kyogenrv_0|krv|id_pc[28]~q ;
wire \kyogenrv_0|krv|id_pc[29]~q ;
wire \kyogenrv_0|krv|id_pc[30]~q ;
wire \kyogenrv_0|krv|id_pc[31]~q ;
wire \pio_0|data_out[0]~q ;
wire \pio_0|data_out[1]~q ;
wire \pio_0|data_out[2]~q ;
wire \pio_0|data_out[3]~q ;
wire \pio_0|data_out[4]~q ;
wire \pio_0|data_out[5]~q ;
wire \pio_0|data_out[6]~q ;
wire \pio_0|data_out[7]~q ;
wire \pio_0|data_out[8]~q ;
wire \pio_0|data_out[9]~q ;
wire \pio_0|data_out[10]~q ;
wire \pio_0|data_out[11]~q ;
wire \pio_0|data_out[12]~q ;
wire \pio_0|data_out[13]~q ;
wire \pio_0|data_out[14]~q ;
wire \pio_0|data_out[15]~q ;
wire \pio_0|data_out[24]~q ;
wire \pio_0|data_out[25]~q ;
wire \pio_0|data_out[26]~q ;
wire \pio_0|data_out[27]~q ;
wire \pio_0|data_out[28]~q ;
wire \pio_0|data_out[29]~q ;
wire \pio_0|data_out[30]~q ;
wire \pio_0|data_out[31]~q ;
wire \kyogenrv_0|krv|mem_alu_out[1]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[1]~q ;
wire \kyogenrv_0|krv|mem_alu_out[0]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[0]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|waitrequest_reset_override~q ;
wire \mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[0]~q ;
wire \kyogenrv_0|krv|mem_ctrl_mem_wr.10~q ;
wire \mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_1|onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ;
wire \rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \kyogenrv_0|krv|mem_rs_1[0]~q ;
wire \kyogenrv_0|krv|Equal68~0_combout ;
wire \kyogenrv_0|krv|Equal73~0_combout ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[0]~16_combout ;
wire \kyogenrv_0|krv|mem_alu_out[2]~q ;
wire \kyogenrv_0|krv|mem_alu_out[3]~q ;
wire \kyogenrv_0|krv|mem_rs_1[1]~q ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[1]~17_combout ;
wire \kyogenrv_0|krv|mem_rs_1[2]~q ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[2]~18_combout ;
wire \kyogenrv_0|krv|mem_rs_1[3]~q ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[3]~19_combout ;
wire \kyogenrv_0|krv|mem_rs_1[4]~q ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[4]~20_combout ;
wire \kyogenrv_0|krv|mem_rs_1[5]~q ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[5]~21_combout ;
wire \kyogenrv_0|krv|mem_rs_1[6]~q ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[6]~22_combout ;
wire \kyogenrv_0|krv|mem_rs_1[7]~q ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[7]~23_combout ;
wire \kyogenrv_0|krv|mem_rs_1[8]~q ;
wire \pio_0|data_out[12]~9_combout ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[8]~24_combout ;
wire \kyogenrv_0|krv|mem_rs_1[9]~q ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[9]~25_combout ;
wire \kyogenrv_0|krv|mem_rs_1[10]~q ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[10]~26_combout ;
wire \kyogenrv_0|krv|mem_rs_1[11]~q ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[11]~27_combout ;
wire \kyogenrv_0|krv|mem_rs_1[12]~q ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[12]~28_combout ;
wire \kyogenrv_0|krv|mem_rs_1[13]~q ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[13]~29_combout ;
wire \kyogenrv_0|krv|mem_rs_1[14]~q ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[14]~30_combout ;
wire \kyogenrv_0|krv|mem_rs_1[15]~q ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[15]~31_combout ;
wire \kyogenrv_0|krv|mem_rs_1[16]~q ;
wire \pio_0|data_out[17]~11_combout ;
wire \kyogenrv_0|krv|mem_rs_1[17]~q ;
wire \kyogenrv_0|krv|mem_rs_1[18]~q ;
wire \kyogenrv_0|krv|mem_rs_1[19]~q ;
wire \kyogenrv_0|krv|mem_rs_1[20]~q ;
wire \kyogenrv_0|krv|mem_rs_1[21]~q ;
wire \kyogenrv_0|krv|mem_rs_1[22]~q ;
wire \kyogenrv_0|krv|mem_rs_1[23]~q ;
wire \pio_0|data_out[27]~13_combout ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[28]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[29]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[30]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[31]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[8]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[9]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[10]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[11]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[12]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[13]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[14]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[15]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[16]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[17]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[18]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[19]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[4]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[3]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[5]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[6]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[7]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[20]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[21]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[22]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[23]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[24]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[25]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[26]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[27]~q ;
wire \pio_0|readdata[1]~combout ;
wire \pio_0|readdata[0]~combout ;
wire \kyogenrv_0|krv|mem_ctrl_mem_wr.00~q ;
wire \kyogenrv_0|krv|w_req~q ;
wire \kyogenrv_0|krv|mem_ctrl_mem_wr.01~q ;
wire \pio_0|readdata[28]~combout ;
wire \pio_0|readdata[29]~combout ;
wire \pio_0|readdata[30]~combout ;
wire \pio_0|readdata[31]~combout ;
wire \pio_0|readdata[8]~combout ;
wire \pio_0|readdata[9]~combout ;
wire \pio_0|readdata[10]~combout ;
wire \pio_0|readdata[11]~combout ;
wire \pio_0|readdata[12]~combout ;
wire \pio_0|readdata[13]~combout ;
wire \pio_0|readdata[14]~combout ;
wire \pio_0|readdata[15]~combout ;
wire \pio_0|readdata[16]~combout ;
wire \pio_0|readdata[17]~combout ;
wire \pio_0|readdata[18]~combout ;
wire \pio_0|readdata[19]~combout ;
wire \pio_0|readdata[4]~combout ;
wire \pio_0|readdata[2]~combout ;
wire \pio_0|readdata[3]~combout ;
wire \pio_0|readdata[5]~combout ;
wire \pio_0|readdata[6]~combout ;
wire \pio_0|readdata[7]~combout ;
wire \pio_0|readdata[20]~combout ;
wire \pio_0|readdata[21]~combout ;
wire \pio_0|readdata[22]~combout ;
wire \pio_0|readdata[23]~combout ;
wire \pio_0|readdata[24]~combout ;
wire \pio_0|readdata[25]~combout ;
wire \pio_0|readdata[26]~combout ;
wire \pio_0|readdata[27]~combout ;
wire \kyogenrv_0|krv|io_imem_add_addr[2]~0_combout ;
wire \kyogenrv_0|krv|io_imem_add_addr[3]~1_combout ;
wire \kyogenrv_0|krv|io_imem_add_addr[4]~2_combout ;
wire \kyogenrv_0|krv|io_imem_add_addr[5]~3_combout ;
wire \kyogenrv_0|krv|io_imem_add_addr[6]~4_combout ;
wire \kyogenrv_0|krv|io_imem_add_addr[7]~5_combout ;
wire \kyogenrv_0|krv|io_imem_add_addr[8]~6_combout ;
wire \kyogenrv_0|krv|io_imem_add_addr[9]~7_combout ;
wire \kyogenrv_0|krv|io_imem_add_addr[10]~8_combout ;
wire \kyogenrv_0|krv|io_imem_add_addr[11]~9_combout ;
wire \kyogenrv_0|krv|io_imem_add_addr[12]~10_combout ;
wire \kyogenrv_0|krv|io_imem_add_addr[13]~11_combout ;
wire \kyogenrv_0|krv|io_imem_add_addr[14]~12_combout ;
wire \mm_interconnect_0|pio_0_s1_translator|read_latency_shift_reg[0]~q ;
wire \kyogenrv_0|krv|_GEN_73[0]~2_combout ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[24]~48_combout ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[25]~49_combout ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[26]~50_combout ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[27]~51_combout ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[28]~52_combout ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[29]~53_combout ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[30]~54_combout ;
wire \kyogenrv_0|krv|io_w_dmem_dat_data[31]~55_combout ;
wire \~GND~combout ;
wire \clk_clk~input_o ;
wire \reset_reset_n~input_o ;


kyogenrv_fpga_altera_reset_controller rst_controller(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

kyogenrv_fpga_kyogenrv_fpga_mm_interconnect_1 mm_interconnect_1(
	.waitrequest_reset_override(\mm_interconnect_0|pio_0_s1_translator|waitrequest_reset_override~q ),
	.read_latency_shift_reg_0(\mm_interconnect_1|onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.w_req(\kyogenrv_0|krv|w_req~q ),
	.clk_clk(\clk_clk~input_o ));

kyogenrv_fpga_kyogenrv_fpga_mm_interconnect_0 mm_interconnect_0(
	.av_readdata_pre_1(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_0(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[0]~q ),
	.waitrequest_reset_override(\mm_interconnect_0|pio_0_s1_translator|waitrequest_reset_override~q ),
	.wait_latency_counter_0(\mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[0]~q ),
	.mem_ctrl_mem_wr10(\kyogenrv_0|krv|mem_ctrl_mem_wr.10~q ),
	.wait_latency_counter_1(\mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[1]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.av_readdata_pre_28(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_29(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_30(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_31(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[31]~q ),
	.av_readdata_pre_8(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_11(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_16(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_17(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_18(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_19(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_4(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_2(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_5(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_20(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_21(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_22(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_23(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_24(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_26(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_27(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[27]~q ),
	.readdata_1(\pio_0|readdata[1]~combout ),
	.readdata_0(\pio_0|readdata[0]~combout ),
	.mem_ctrl_mem_wr00(\kyogenrv_0|krv|mem_ctrl_mem_wr.00~q ),
	.mem_ctrl_mem_wr01(\kyogenrv_0|krv|mem_ctrl_mem_wr.01~q ),
	.readdata_28(\pio_0|readdata[28]~combout ),
	.readdata_29(\pio_0|readdata[29]~combout ),
	.readdata_30(\pio_0|readdata[30]~combout ),
	.readdata_31(\pio_0|readdata[31]~combout ),
	.readdata_8(\pio_0|readdata[8]~combout ),
	.readdata_9(\pio_0|readdata[9]~combout ),
	.readdata_10(\pio_0|readdata[10]~combout ),
	.readdata_11(\pio_0|readdata[11]~combout ),
	.readdata_12(\pio_0|readdata[12]~combout ),
	.readdata_13(\pio_0|readdata[13]~combout ),
	.readdata_14(\pio_0|readdata[14]~combout ),
	.readdata_15(\pio_0|readdata[15]~combout ),
	.readdata_16(\pio_0|readdata[16]~combout ),
	.readdata_17(\pio_0|readdata[17]~combout ),
	.readdata_18(\pio_0|readdata[18]~combout ),
	.readdata_19(\pio_0|readdata[19]~combout ),
	.readdata_4(\pio_0|readdata[4]~combout ),
	.readdata_2(\pio_0|readdata[2]~combout ),
	.readdata_3(\pio_0|readdata[3]~combout ),
	.readdata_5(\pio_0|readdata[5]~combout ),
	.readdata_6(\pio_0|readdata[6]~combout ),
	.readdata_7(\pio_0|readdata[7]~combout ),
	.readdata_20(\pio_0|readdata[20]~combout ),
	.readdata_21(\pio_0|readdata[21]~combout ),
	.readdata_22(\pio_0|readdata[22]~combout ),
	.readdata_23(\pio_0|readdata[23]~combout ),
	.readdata_24(\pio_0|readdata[24]~combout ),
	.readdata_25(\pio_0|readdata[25]~combout ),
	.readdata_26(\pio_0|readdata[26]~combout ),
	.readdata_27(\pio_0|readdata[27]~combout ),
	.read_latency_shift_reg_0(\mm_interconnect_0|pio_0_s1_translator|read_latency_shift_reg[0]~q ),
	.clk_clk(\clk_clk~input_o ));

kyogenrv_fpga_kyogenrv_fpga_pio_0 pio_0(
	.data_out_16(\pio_0|data_out[16]~q ),
	.data_out_17(\pio_0|data_out[17]~q ),
	.data_out_18(\pio_0|data_out[18]~q ),
	.data_out_19(\pio_0|data_out[19]~q ),
	.data_out_20(\pio_0|data_out[20]~q ),
	.data_out_21(\pio_0|data_out[21]~q ),
	.data_out_22(\pio_0|data_out[22]~q ),
	.data_out_23(\pio_0|data_out[23]~q ),
	.data_out_0(\pio_0|data_out[0]~q ),
	.data_out_1(\pio_0|data_out[1]~q ),
	.data_out_2(\pio_0|data_out[2]~q ),
	.data_out_3(\pio_0|data_out[3]~q ),
	.data_out_4(\pio_0|data_out[4]~q ),
	.data_out_5(\pio_0|data_out[5]~q ),
	.data_out_6(\pio_0|data_out[6]~q ),
	.data_out_7(\pio_0|data_out[7]~q ),
	.data_out_8(\pio_0|data_out[8]~q ),
	.data_out_9(\pio_0|data_out[9]~q ),
	.data_out_10(\pio_0|data_out[10]~q ),
	.data_out_11(\pio_0|data_out[11]~q ),
	.data_out_12(\pio_0|data_out[12]~q ),
	.data_out_13(\pio_0|data_out[13]~q ),
	.data_out_14(\pio_0|data_out[14]~q ),
	.data_out_15(\pio_0|data_out[15]~q ),
	.data_out_24(\pio_0|data_out[24]~q ),
	.data_out_25(\pio_0|data_out[25]~q ),
	.data_out_26(\pio_0|data_out[26]~q ),
	.data_out_27(\pio_0|data_out[27]~q ),
	.data_out_28(\pio_0|data_out[28]~q ),
	.data_out_29(\pio_0|data_out[29]~q ),
	.data_out_30(\pio_0|data_out[30]~q ),
	.data_out_31(\pio_0|data_out[31]~q ),
	.mem_alu_out_1(\kyogenrv_0|krv|mem_alu_out[1]~q ),
	.mem_alu_out_0(\kyogenrv_0|krv|mem_alu_out[0]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[0]~q ),
	.mem_ctrl_mem_wr10(\kyogenrv_0|krv|mem_ctrl_mem_wr.10~q ),
	.wait_latency_counter_1(\mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[1]~q ),
	.reset_n(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.mem_rs_1_0(\kyogenrv_0|krv|mem_rs_1[0]~q ),
	.Equal68(\kyogenrv_0|krv|Equal68~0_combout ),
	.Equal73(\kyogenrv_0|krv|Equal73~0_combout ),
	.writedata({\kyogenrv_0|krv|io_w_dmem_dat_data[31]~55_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[30]~54_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[29]~53_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[28]~52_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[27]~51_combout ,
\kyogenrv_0|krv|io_w_dmem_dat_data[26]~50_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[25]~49_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[24]~48_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\kyogenrv_0|krv|io_w_dmem_dat_data[15]~31_combout ,
\kyogenrv_0|krv|io_w_dmem_dat_data[14]~30_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[13]~29_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[12]~28_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[11]~27_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[10]~26_combout ,
\kyogenrv_0|krv|io_w_dmem_dat_data[9]~25_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[8]~24_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[7]~23_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[6]~22_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[5]~21_combout ,
\kyogenrv_0|krv|io_w_dmem_dat_data[4]~20_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[3]~19_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[2]~18_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[1]~17_combout ,\kyogenrv_0|krv|io_w_dmem_dat_data[0]~16_combout }),
	.mem_alu_out_2(\kyogenrv_0|krv|mem_alu_out[2]~q ),
	.mem_alu_out_3(\kyogenrv_0|krv|mem_alu_out[3]~q ),
	.mem_rs_1_1(\kyogenrv_0|krv|mem_rs_1[1]~q ),
	.mem_rs_1_2(\kyogenrv_0|krv|mem_rs_1[2]~q ),
	.mem_rs_1_3(\kyogenrv_0|krv|mem_rs_1[3]~q ),
	.mem_rs_1_4(\kyogenrv_0|krv|mem_rs_1[4]~q ),
	.mem_rs_1_5(\kyogenrv_0|krv|mem_rs_1[5]~q ),
	.mem_rs_1_6(\kyogenrv_0|krv|mem_rs_1[6]~q ),
	.mem_rs_1_7(\kyogenrv_0|krv|mem_rs_1[7]~q ),
	.mem_rs_1_8(\kyogenrv_0|krv|mem_rs_1[8]~q ),
	.data_out_121(\pio_0|data_out[12]~9_combout ),
	.mem_rs_1_9(\kyogenrv_0|krv|mem_rs_1[9]~q ),
	.mem_rs_1_10(\kyogenrv_0|krv|mem_rs_1[10]~q ),
	.mem_rs_1_11(\kyogenrv_0|krv|mem_rs_1[11]~q ),
	.mem_rs_1_12(\kyogenrv_0|krv|mem_rs_1[12]~q ),
	.mem_rs_1_13(\kyogenrv_0|krv|mem_rs_1[13]~q ),
	.mem_rs_1_14(\kyogenrv_0|krv|mem_rs_1[14]~q ),
	.mem_rs_1_15(\kyogenrv_0|krv|mem_rs_1[15]~q ),
	.mem_rs_1_16(\kyogenrv_0|krv|mem_rs_1[16]~q ),
	.data_out_171(\pio_0|data_out[17]~11_combout ),
	.mem_rs_1_17(\kyogenrv_0|krv|mem_rs_1[17]~q ),
	.mem_rs_1_18(\kyogenrv_0|krv|mem_rs_1[18]~q ),
	.mem_rs_1_19(\kyogenrv_0|krv|mem_rs_1[19]~q ),
	.mem_rs_1_20(\kyogenrv_0|krv|mem_rs_1[20]~q ),
	.mem_rs_1_21(\kyogenrv_0|krv|mem_rs_1[21]~q ),
	.mem_rs_1_22(\kyogenrv_0|krv|mem_rs_1[22]~q ),
	.mem_rs_1_23(\kyogenrv_0|krv|mem_rs_1[23]~q ),
	.data_out_271(\pio_0|data_out[27]~13_combout ),
	.readdata_1(\pio_0|readdata[1]~combout ),
	.readdata_0(\pio_0|readdata[0]~combout ),
	.readdata_28(\pio_0|readdata[28]~combout ),
	.readdata_29(\pio_0|readdata[29]~combout ),
	.readdata_30(\pio_0|readdata[30]~combout ),
	.readdata_31(\pio_0|readdata[31]~combout ),
	.readdata_8(\pio_0|readdata[8]~combout ),
	.readdata_9(\pio_0|readdata[9]~combout ),
	.readdata_10(\pio_0|readdata[10]~combout ),
	.readdata_11(\pio_0|readdata[11]~combout ),
	.readdata_12(\pio_0|readdata[12]~combout ),
	.readdata_13(\pio_0|readdata[13]~combout ),
	.readdata_14(\pio_0|readdata[14]~combout ),
	.readdata_15(\pio_0|readdata[15]~combout ),
	.readdata_16(\pio_0|readdata[16]~combout ),
	.readdata_17(\pio_0|readdata[17]~combout ),
	.readdata_18(\pio_0|readdata[18]~combout ),
	.readdata_19(\pio_0|readdata[19]~combout ),
	.readdata_4(\pio_0|readdata[4]~combout ),
	.readdata_2(\pio_0|readdata[2]~combout ),
	.readdata_3(\pio_0|readdata[3]~combout ),
	.readdata_5(\pio_0|readdata[5]~combout ),
	.readdata_6(\pio_0|readdata[6]~combout ),
	.readdata_7(\pio_0|readdata[7]~combout ),
	.readdata_20(\pio_0|readdata[20]~combout ),
	.readdata_21(\pio_0|readdata[21]~combout ),
	.readdata_22(\pio_0|readdata[22]~combout ),
	.readdata_23(\pio_0|readdata[23]~combout ),
	.readdata_24(\pio_0|readdata[24]~combout ),
	.readdata_25(\pio_0|readdata[25]~combout ),
	.readdata_26(\pio_0|readdata[26]~combout ),
	.readdata_27(\pio_0|readdata[27]~combout ),
	._GEN_73_0(\kyogenrv_0|krv|_GEN_73[0]~2_combout ),
	.clk(\clk_clk~input_o ));

kyogenrv_fpga_kyogenrv_fpga_onchip_memory2_0 onchip_memory2_0(
	.q_a_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_24(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_6(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_7(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_11(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_25(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_30(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_0(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_2(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_26(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_27(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_31(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_28(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_29(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ),
	.w_req(\kyogenrv_0|krv|w_req~q ),
	.io_imem_add_addr_2(\kyogenrv_0|krv|io_imem_add_addr[2]~0_combout ),
	.io_imem_add_addr_3(\kyogenrv_0|krv|io_imem_add_addr[3]~1_combout ),
	.io_imem_add_addr_4(\kyogenrv_0|krv|io_imem_add_addr[4]~2_combout ),
	.io_imem_add_addr_5(\kyogenrv_0|krv|io_imem_add_addr[5]~3_combout ),
	.io_imem_add_addr_6(\kyogenrv_0|krv|io_imem_add_addr[6]~4_combout ),
	.io_imem_add_addr_7(\kyogenrv_0|krv|io_imem_add_addr[7]~5_combout ),
	.io_imem_add_addr_8(\kyogenrv_0|krv|io_imem_add_addr[8]~6_combout ),
	.io_imem_add_addr_9(\kyogenrv_0|krv|io_imem_add_addr[9]~7_combout ),
	.io_imem_add_addr_10(\kyogenrv_0|krv|io_imem_add_addr[10]~8_combout ),
	.io_imem_add_addr_11(\kyogenrv_0|krv|io_imem_add_addr[11]~9_combout ),
	.io_imem_add_addr_12(\kyogenrv_0|krv|io_imem_add_addr[12]~10_combout ),
	.io_imem_add_addr_13(\kyogenrv_0|krv|io_imem_add_addr[13]~11_combout ),
	.io_imem_add_addr_14(\kyogenrv_0|krv|io_imem_add_addr[14]~12_combout ),
	.GND_port(\~GND~combout ),
	.clk_clk(\clk_clk~input_o ));

kyogenrv_fpga_kyogenrv_fpga_avalonMM kyogenrv_0(
	.q_a_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_24(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_6(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_7(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_11(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_25(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_30(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_0(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_2(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_26(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_27(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_31(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_28(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_29(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ),
	.id_npc_0(\kyogenrv_0|krv|id_npc[0]~q ),
	.id_npc_1(\kyogenrv_0|krv|id_npc[1]~q ),
	.id_pc_2(\kyogenrv_0|krv|id_pc[2]~q ),
	.id_pc_3(\kyogenrv_0|krv|id_pc[3]~q ),
	.id_pc_4(\kyogenrv_0|krv|id_pc[4]~q ),
	.id_pc_5(\kyogenrv_0|krv|id_pc[5]~q ),
	.id_pc_6(\kyogenrv_0|krv|id_pc[6]~q ),
	.id_pc_7(\kyogenrv_0|krv|id_pc[7]~q ),
	.id_pc_8(\kyogenrv_0|krv|id_pc[8]~q ),
	.id_pc_9(\kyogenrv_0|krv|id_pc[9]~q ),
	.id_pc_10(\kyogenrv_0|krv|id_pc[10]~q ),
	.id_pc_11(\kyogenrv_0|krv|id_pc[11]~q ),
	.id_pc_12(\kyogenrv_0|krv|id_pc[12]~q ),
	.id_pc_13(\kyogenrv_0|krv|id_pc[13]~q ),
	.id_pc_14(\kyogenrv_0|krv|id_pc[14]~q ),
	.id_pc_15(\kyogenrv_0|krv|id_pc[15]~q ),
	.id_pc_16(\kyogenrv_0|krv|id_pc[16]~q ),
	.id_pc_17(\kyogenrv_0|krv|id_pc[17]~q ),
	.id_pc_18(\kyogenrv_0|krv|id_pc[18]~q ),
	.id_pc_19(\kyogenrv_0|krv|id_pc[19]~q ),
	.id_pc_20(\kyogenrv_0|krv|id_pc[20]~q ),
	.id_pc_21(\kyogenrv_0|krv|id_pc[21]~q ),
	.id_pc_22(\kyogenrv_0|krv|id_pc[22]~q ),
	.id_pc_23(\kyogenrv_0|krv|id_pc[23]~q ),
	.id_pc_24(\kyogenrv_0|krv|id_pc[24]~q ),
	.id_pc_25(\kyogenrv_0|krv|id_pc[25]~q ),
	.id_pc_26(\kyogenrv_0|krv|id_pc[26]~q ),
	.id_pc_27(\kyogenrv_0|krv|id_pc[27]~q ),
	.id_pc_28(\kyogenrv_0|krv|id_pc[28]~q ),
	.id_pc_29(\kyogenrv_0|krv|id_pc[29]~q ),
	.id_pc_30(\kyogenrv_0|krv|id_pc[30]~q ),
	.id_pc_31(\kyogenrv_0|krv|id_pc[31]~q ),
	.mem_alu_out_1(\kyogenrv_0|krv|mem_alu_out[1]~q ),
	.av_readdata_pre_1(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[1]~q ),
	.mem_alu_out_0(\kyogenrv_0|krv|mem_alu_out[0]~q ),
	.av_readdata_pre_0(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[0]~q ),
	.waitrequest_reset_override(\mm_interconnect_0|pio_0_s1_translator|waitrequest_reset_override~q ),
	.wait_latency_counter_0(\mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[0]~q ),
	.mem_ctrl_mem_wr10(\kyogenrv_0|krv|mem_ctrl_mem_wr.10~q ),
	.wait_latency_counter_1(\mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[1]~q ),
	.read_latency_shift_reg_0(\mm_interconnect_1|onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.mem_rs_1_0(\kyogenrv_0|krv|mem_rs_1[0]~q ),
	.Equal68(\kyogenrv_0|krv|Equal68~0_combout ),
	.Equal73(\kyogenrv_0|krv|Equal73~0_combout ),
	.io_w_dmem_dat_data_0(\kyogenrv_0|krv|io_w_dmem_dat_data[0]~16_combout ),
	.mem_alu_out_2(\kyogenrv_0|krv|mem_alu_out[2]~q ),
	.mem_alu_out_3(\kyogenrv_0|krv|mem_alu_out[3]~q ),
	.mem_rs_1_1(\kyogenrv_0|krv|mem_rs_1[1]~q ),
	.io_w_dmem_dat_data_1(\kyogenrv_0|krv|io_w_dmem_dat_data[1]~17_combout ),
	.mem_rs_1_2(\kyogenrv_0|krv|mem_rs_1[2]~q ),
	.io_w_dmem_dat_data_2(\kyogenrv_0|krv|io_w_dmem_dat_data[2]~18_combout ),
	.mem_rs_1_3(\kyogenrv_0|krv|mem_rs_1[3]~q ),
	.io_w_dmem_dat_data_3(\kyogenrv_0|krv|io_w_dmem_dat_data[3]~19_combout ),
	.mem_rs_1_4(\kyogenrv_0|krv|mem_rs_1[4]~q ),
	.io_w_dmem_dat_data_4(\kyogenrv_0|krv|io_w_dmem_dat_data[4]~20_combout ),
	.mem_rs_1_5(\kyogenrv_0|krv|mem_rs_1[5]~q ),
	.io_w_dmem_dat_data_5(\kyogenrv_0|krv|io_w_dmem_dat_data[5]~21_combout ),
	.mem_rs_1_6(\kyogenrv_0|krv|mem_rs_1[6]~q ),
	.io_w_dmem_dat_data_6(\kyogenrv_0|krv|io_w_dmem_dat_data[6]~22_combout ),
	.mem_rs_1_7(\kyogenrv_0|krv|mem_rs_1[7]~q ),
	.io_w_dmem_dat_data_7(\kyogenrv_0|krv|io_w_dmem_dat_data[7]~23_combout ),
	.mem_rs_1_8(\kyogenrv_0|krv|mem_rs_1[8]~q ),
	.data_out_12(\pio_0|data_out[12]~9_combout ),
	.io_w_dmem_dat_data_8(\kyogenrv_0|krv|io_w_dmem_dat_data[8]~24_combout ),
	.mem_rs_1_9(\kyogenrv_0|krv|mem_rs_1[9]~q ),
	.io_w_dmem_dat_data_9(\kyogenrv_0|krv|io_w_dmem_dat_data[9]~25_combout ),
	.mem_rs_1_10(\kyogenrv_0|krv|mem_rs_1[10]~q ),
	.io_w_dmem_dat_data_10(\kyogenrv_0|krv|io_w_dmem_dat_data[10]~26_combout ),
	.mem_rs_1_11(\kyogenrv_0|krv|mem_rs_1[11]~q ),
	.io_w_dmem_dat_data_11(\kyogenrv_0|krv|io_w_dmem_dat_data[11]~27_combout ),
	.mem_rs_1_12(\kyogenrv_0|krv|mem_rs_1[12]~q ),
	.io_w_dmem_dat_data_12(\kyogenrv_0|krv|io_w_dmem_dat_data[12]~28_combout ),
	.mem_rs_1_13(\kyogenrv_0|krv|mem_rs_1[13]~q ),
	.io_w_dmem_dat_data_13(\kyogenrv_0|krv|io_w_dmem_dat_data[13]~29_combout ),
	.mem_rs_1_14(\kyogenrv_0|krv|mem_rs_1[14]~q ),
	.io_w_dmem_dat_data_14(\kyogenrv_0|krv|io_w_dmem_dat_data[14]~30_combout ),
	.mem_rs_1_15(\kyogenrv_0|krv|mem_rs_1[15]~q ),
	.io_w_dmem_dat_data_15(\kyogenrv_0|krv|io_w_dmem_dat_data[15]~31_combout ),
	.mem_rs_1_16(\kyogenrv_0|krv|mem_rs_1[16]~q ),
	.data_out_17(\pio_0|data_out[17]~11_combout ),
	.mem_rs_1_17(\kyogenrv_0|krv|mem_rs_1[17]~q ),
	.mem_rs_1_18(\kyogenrv_0|krv|mem_rs_1[18]~q ),
	.mem_rs_1_19(\kyogenrv_0|krv|mem_rs_1[19]~q ),
	.mem_rs_1_20(\kyogenrv_0|krv|mem_rs_1[20]~q ),
	.mem_rs_1_21(\kyogenrv_0|krv|mem_rs_1[21]~q ),
	.mem_rs_1_22(\kyogenrv_0|krv|mem_rs_1[22]~q ),
	.mem_rs_1_23(\kyogenrv_0|krv|mem_rs_1[23]~q ),
	.data_out_27(\pio_0|data_out[27]~13_combout ),
	.av_readdata_pre_28(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_29(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_30(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_31(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[31]~q ),
	.av_readdata_pre_8(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_11(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_16(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_17(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_18(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_19(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_4(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_2(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_5(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_20(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_21(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_22(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_23(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_24(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_26(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_27(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[27]~q ),
	.mem_ctrl_mem_wr00(\kyogenrv_0|krv|mem_ctrl_mem_wr.00~q ),
	.w_req(\kyogenrv_0|krv|w_req~q ),
	.mem_ctrl_mem_wr01(\kyogenrv_0|krv|mem_ctrl_mem_wr.01~q ),
	.io_imem_add_addr_2(\kyogenrv_0|krv|io_imem_add_addr[2]~0_combout ),
	.io_imem_add_addr_3(\kyogenrv_0|krv|io_imem_add_addr[3]~1_combout ),
	.io_imem_add_addr_4(\kyogenrv_0|krv|io_imem_add_addr[4]~2_combout ),
	.io_imem_add_addr_5(\kyogenrv_0|krv|io_imem_add_addr[5]~3_combout ),
	.io_imem_add_addr_6(\kyogenrv_0|krv|io_imem_add_addr[6]~4_combout ),
	.io_imem_add_addr_7(\kyogenrv_0|krv|io_imem_add_addr[7]~5_combout ),
	.io_imem_add_addr_8(\kyogenrv_0|krv|io_imem_add_addr[8]~6_combout ),
	.io_imem_add_addr_9(\kyogenrv_0|krv|io_imem_add_addr[9]~7_combout ),
	.io_imem_add_addr_10(\kyogenrv_0|krv|io_imem_add_addr[10]~8_combout ),
	.io_imem_add_addr_11(\kyogenrv_0|krv|io_imem_add_addr[11]~9_combout ),
	.io_imem_add_addr_12(\kyogenrv_0|krv|io_imem_add_addr[12]~10_combout ),
	.io_imem_add_addr_13(\kyogenrv_0|krv|io_imem_add_addr[13]~11_combout ),
	.io_imem_add_addr_14(\kyogenrv_0|krv|io_imem_add_addr[14]~12_combout ),
	.read_latency_shift_reg_01(\mm_interconnect_0|pio_0_s1_translator|read_latency_shift_reg[0]~q ),
	._GEN_73_0(\kyogenrv_0|krv|_GEN_73[0]~2_combout ),
	.io_w_dmem_dat_data_24(\kyogenrv_0|krv|io_w_dmem_dat_data[24]~48_combout ),
	.io_w_dmem_dat_data_25(\kyogenrv_0|krv|io_w_dmem_dat_data[25]~49_combout ),
	.io_w_dmem_dat_data_26(\kyogenrv_0|krv|io_w_dmem_dat_data[26]~50_combout ),
	.io_w_dmem_dat_data_27(\kyogenrv_0|krv|io_w_dmem_dat_data[27]~51_combout ),
	.io_w_dmem_dat_data_28(\kyogenrv_0|krv|io_w_dmem_dat_data[28]~52_combout ),
	.io_w_dmem_dat_data_29(\kyogenrv_0|krv|io_w_dmem_dat_data[29]~53_combout ),
	.io_w_dmem_dat_data_30(\kyogenrv_0|krv|io_w_dmem_dat_data[30]~54_combout ),
	.io_w_dmem_dat_data_31(\kyogenrv_0|krv|io_w_dmem_dat_data[31]~55_combout ),
	.clk_clk(\clk_clk~input_o ));

cyclone10lp_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

assign \clk_clk~input_o  = clk_clk;

assign \reset_reset_n~input_o  = reset_reset_n;

assign kyogenrv_0_counter_readdata[0] = \kyogenrv_0|krv|id_npc[0]~q ;

assign kyogenrv_0_counter_readdata[1] = \kyogenrv_0|krv|id_npc[1]~q ;

assign kyogenrv_0_counter_readdata[2] = \kyogenrv_0|krv|id_pc[2]~q ;

assign kyogenrv_0_counter_readdata[3] = \kyogenrv_0|krv|id_pc[3]~q ;

assign kyogenrv_0_counter_readdata[4] = \kyogenrv_0|krv|id_pc[4]~q ;

assign kyogenrv_0_counter_readdata[5] = \kyogenrv_0|krv|id_pc[5]~q ;

assign kyogenrv_0_counter_readdata[6] = \kyogenrv_0|krv|id_pc[6]~q ;

assign kyogenrv_0_counter_readdata[7] = \kyogenrv_0|krv|id_pc[7]~q ;

assign kyogenrv_0_counter_readdata[8] = \kyogenrv_0|krv|id_pc[8]~q ;

assign kyogenrv_0_counter_readdata[9] = \kyogenrv_0|krv|id_pc[9]~q ;

assign kyogenrv_0_counter_readdata[10] = \kyogenrv_0|krv|id_pc[10]~q ;

assign kyogenrv_0_counter_readdata[11] = \kyogenrv_0|krv|id_pc[11]~q ;

assign kyogenrv_0_counter_readdata[12] = \kyogenrv_0|krv|id_pc[12]~q ;

assign kyogenrv_0_counter_readdata[13] = \kyogenrv_0|krv|id_pc[13]~q ;

assign kyogenrv_0_counter_readdata[14] = \kyogenrv_0|krv|id_pc[14]~q ;

assign kyogenrv_0_counter_readdata[15] = \kyogenrv_0|krv|id_pc[15]~q ;

assign kyogenrv_0_counter_readdata[16] = \kyogenrv_0|krv|id_pc[16]~q ;

assign kyogenrv_0_counter_readdata[17] = \kyogenrv_0|krv|id_pc[17]~q ;

assign kyogenrv_0_counter_readdata[18] = \kyogenrv_0|krv|id_pc[18]~q ;

assign kyogenrv_0_counter_readdata[19] = \kyogenrv_0|krv|id_pc[19]~q ;

assign kyogenrv_0_counter_readdata[20] = \kyogenrv_0|krv|id_pc[20]~q ;

assign kyogenrv_0_counter_readdata[21] = \kyogenrv_0|krv|id_pc[21]~q ;

assign kyogenrv_0_counter_readdata[22] = \kyogenrv_0|krv|id_pc[22]~q ;

assign kyogenrv_0_counter_readdata[23] = \kyogenrv_0|krv|id_pc[23]~q ;

assign kyogenrv_0_counter_readdata[24] = \kyogenrv_0|krv|id_pc[24]~q ;

assign kyogenrv_0_counter_readdata[25] = \kyogenrv_0|krv|id_pc[25]~q ;

assign kyogenrv_0_counter_readdata[26] = \kyogenrv_0|krv|id_pc[26]~q ;

assign kyogenrv_0_counter_readdata[27] = \kyogenrv_0|krv|id_pc[27]~q ;

assign kyogenrv_0_counter_readdata[28] = \kyogenrv_0|krv|id_pc[28]~q ;

assign kyogenrv_0_counter_readdata[29] = \kyogenrv_0|krv|id_pc[29]~q ;

assign kyogenrv_0_counter_readdata[30] = \kyogenrv_0|krv|id_pc[30]~q ;

assign kyogenrv_0_counter_readdata[31] = \kyogenrv_0|krv|id_pc[31]~q ;

assign pio_0_external_connection_export[0] = \pio_0|data_out[0]~q ;

assign pio_0_external_connection_export[1] = \pio_0|data_out[1]~q ;

assign pio_0_external_connection_export[2] = \pio_0|data_out[2]~q ;

assign pio_0_external_connection_export[3] = \pio_0|data_out[3]~q ;

assign pio_0_external_connection_export[4] = \pio_0|data_out[4]~q ;

assign pio_0_external_connection_export[5] = \pio_0|data_out[5]~q ;

assign pio_0_external_connection_export[6] = \pio_0|data_out[6]~q ;

assign pio_0_external_connection_export[7] = \pio_0|data_out[7]~q ;

assign pio_0_external_connection_export[8] = \pio_0|data_out[8]~q ;

assign pio_0_external_connection_export[9] = \pio_0|data_out[9]~q ;

assign pio_0_external_connection_export[10] = \pio_0|data_out[10]~q ;

assign pio_0_external_connection_export[11] = \pio_0|data_out[11]~q ;

assign pio_0_external_connection_export[12] = \pio_0|data_out[12]~q ;

assign pio_0_external_connection_export[13] = \pio_0|data_out[13]~q ;

assign pio_0_external_connection_export[14] = \pio_0|data_out[14]~q ;

assign pio_0_external_connection_export[15] = \pio_0|data_out[15]~q ;

assign pio_0_external_connection_export[16] = \pio_0|data_out[16]~q ;

assign pio_0_external_connection_export[17] = \pio_0|data_out[17]~q ;

assign pio_0_external_connection_export[18] = \pio_0|data_out[18]~q ;

assign pio_0_external_connection_export[19] = \pio_0|data_out[19]~q ;

assign pio_0_external_connection_export[20] = \pio_0|data_out[20]~q ;

assign pio_0_external_connection_export[21] = \pio_0|data_out[21]~q ;

assign pio_0_external_connection_export[22] = \pio_0|data_out[22]~q ;

assign pio_0_external_connection_export[23] = \pio_0|data_out[23]~q ;

assign pio_0_external_connection_export[24] = \pio_0|data_out[24]~q ;

assign pio_0_external_connection_export[25] = \pio_0|data_out[25]~q ;

assign pio_0_external_connection_export[26] = \pio_0|data_out[26]~q ;

assign pio_0_external_connection_export[27] = \pio_0|data_out[27]~q ;

assign pio_0_external_connection_export[28] = \pio_0|data_out[28]~q ;

assign pio_0_external_connection_export[29] = \pio_0|data_out[29]~q ;

assign pio_0_external_connection_export[30] = \pio_0|data_out[30]~q ;

assign pio_0_external_connection_export[31] = \pio_0|data_out[31]~q ;

endmodule

module kyogenrv_fpga_altera_reset_controller (
	altera_reset_synchronizer_int_chain_out,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



kyogenrv_fpga_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

endmodule

module kyogenrv_fpga_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module kyogenrv_fpga_kyogenrv_fpga_avalonMM (
	q_a_16,
	q_a_15,
	q_a_18,
	q_a_17,
	q_a_19,
	q_a_21,
	q_a_20,
	q_a_23,
	q_a_22,
	q_a_24,
	q_a_14,
	q_a_13,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	q_a_12,
	q_a_10,
	q_a_11,
	q_a_25,
	q_a_30,
	q_a_0,
	q_a_1,
	q_a_3,
	q_a_2,
	q_a_4,
	q_a_26,
	q_a_27,
	q_a_31,
	q_a_28,
	q_a_29,
	id_npc_0,
	id_npc_1,
	id_pc_2,
	id_pc_3,
	id_pc_4,
	id_pc_5,
	id_pc_6,
	id_pc_7,
	id_pc_8,
	id_pc_9,
	id_pc_10,
	id_pc_11,
	id_pc_12,
	id_pc_13,
	id_pc_14,
	id_pc_15,
	id_pc_16,
	id_pc_17,
	id_pc_18,
	id_pc_19,
	id_pc_20,
	id_pc_21,
	id_pc_22,
	id_pc_23,
	id_pc_24,
	id_pc_25,
	id_pc_26,
	id_pc_27,
	id_pc_28,
	id_pc_29,
	id_pc_30,
	id_pc_31,
	mem_alu_out_1,
	av_readdata_pre_1,
	mem_alu_out_0,
	av_readdata_pre_0,
	waitrequest_reset_override,
	wait_latency_counter_0,
	mem_ctrl_mem_wr10,
	wait_latency_counter_1,
	read_latency_shift_reg_0,
	altera_reset_synchronizer_int_chain_out,
	mem_rs_1_0,
	Equal68,
	Equal73,
	io_w_dmem_dat_data_0,
	mem_alu_out_2,
	mem_alu_out_3,
	mem_rs_1_1,
	io_w_dmem_dat_data_1,
	mem_rs_1_2,
	io_w_dmem_dat_data_2,
	mem_rs_1_3,
	io_w_dmem_dat_data_3,
	mem_rs_1_4,
	io_w_dmem_dat_data_4,
	mem_rs_1_5,
	io_w_dmem_dat_data_5,
	mem_rs_1_6,
	io_w_dmem_dat_data_6,
	mem_rs_1_7,
	io_w_dmem_dat_data_7,
	mem_rs_1_8,
	data_out_12,
	io_w_dmem_dat_data_8,
	mem_rs_1_9,
	io_w_dmem_dat_data_9,
	mem_rs_1_10,
	io_w_dmem_dat_data_10,
	mem_rs_1_11,
	io_w_dmem_dat_data_11,
	mem_rs_1_12,
	io_w_dmem_dat_data_12,
	mem_rs_1_13,
	io_w_dmem_dat_data_13,
	mem_rs_1_14,
	io_w_dmem_dat_data_14,
	mem_rs_1_15,
	io_w_dmem_dat_data_15,
	mem_rs_1_16,
	data_out_17,
	mem_rs_1_17,
	mem_rs_1_18,
	mem_rs_1_19,
	mem_rs_1_20,
	mem_rs_1_21,
	mem_rs_1_22,
	mem_rs_1_23,
	data_out_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_30,
	av_readdata_pre_31,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata_pre_18,
	av_readdata_pre_19,
	av_readdata_pre_4,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_20,
	av_readdata_pre_21,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_27,
	mem_ctrl_mem_wr00,
	w_req,
	mem_ctrl_mem_wr01,
	io_imem_add_addr_2,
	io_imem_add_addr_3,
	io_imem_add_addr_4,
	io_imem_add_addr_5,
	io_imem_add_addr_6,
	io_imem_add_addr_7,
	io_imem_add_addr_8,
	io_imem_add_addr_9,
	io_imem_add_addr_10,
	io_imem_add_addr_11,
	io_imem_add_addr_12,
	io_imem_add_addr_13,
	io_imem_add_addr_14,
	read_latency_shift_reg_01,
	_GEN_73_0,
	io_w_dmem_dat_data_24,
	io_w_dmem_dat_data_25,
	io_w_dmem_dat_data_26,
	io_w_dmem_dat_data_27,
	io_w_dmem_dat_data_28,
	io_w_dmem_dat_data_29,
	io_w_dmem_dat_data_30,
	io_w_dmem_dat_data_31,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	q_a_16;
input 	q_a_15;
input 	q_a_18;
input 	q_a_17;
input 	q_a_19;
input 	q_a_21;
input 	q_a_20;
input 	q_a_23;
input 	q_a_22;
input 	q_a_24;
input 	q_a_14;
input 	q_a_13;
input 	q_a_5;
input 	q_a_6;
input 	q_a_7;
input 	q_a_8;
input 	q_a_9;
input 	q_a_12;
input 	q_a_10;
input 	q_a_11;
input 	q_a_25;
input 	q_a_30;
input 	q_a_0;
input 	q_a_1;
input 	q_a_3;
input 	q_a_2;
input 	q_a_4;
input 	q_a_26;
input 	q_a_27;
input 	q_a_31;
input 	q_a_28;
input 	q_a_29;
output 	id_npc_0;
output 	id_npc_1;
output 	id_pc_2;
output 	id_pc_3;
output 	id_pc_4;
output 	id_pc_5;
output 	id_pc_6;
output 	id_pc_7;
output 	id_pc_8;
output 	id_pc_9;
output 	id_pc_10;
output 	id_pc_11;
output 	id_pc_12;
output 	id_pc_13;
output 	id_pc_14;
output 	id_pc_15;
output 	id_pc_16;
output 	id_pc_17;
output 	id_pc_18;
output 	id_pc_19;
output 	id_pc_20;
output 	id_pc_21;
output 	id_pc_22;
output 	id_pc_23;
output 	id_pc_24;
output 	id_pc_25;
output 	id_pc_26;
output 	id_pc_27;
output 	id_pc_28;
output 	id_pc_29;
output 	id_pc_30;
output 	id_pc_31;
output 	mem_alu_out_1;
input 	av_readdata_pre_1;
output 	mem_alu_out_0;
input 	av_readdata_pre_0;
input 	waitrequest_reset_override;
input 	wait_latency_counter_0;
output 	mem_ctrl_mem_wr10;
input 	wait_latency_counter_1;
input 	read_latency_shift_reg_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	mem_rs_1_0;
output 	Equal68;
output 	Equal73;
output 	io_w_dmem_dat_data_0;
output 	mem_alu_out_2;
output 	mem_alu_out_3;
output 	mem_rs_1_1;
output 	io_w_dmem_dat_data_1;
output 	mem_rs_1_2;
output 	io_w_dmem_dat_data_2;
output 	mem_rs_1_3;
output 	io_w_dmem_dat_data_3;
output 	mem_rs_1_4;
output 	io_w_dmem_dat_data_4;
output 	mem_rs_1_5;
output 	io_w_dmem_dat_data_5;
output 	mem_rs_1_6;
output 	io_w_dmem_dat_data_6;
output 	mem_rs_1_7;
output 	io_w_dmem_dat_data_7;
output 	mem_rs_1_8;
input 	data_out_12;
output 	io_w_dmem_dat_data_8;
output 	mem_rs_1_9;
output 	io_w_dmem_dat_data_9;
output 	mem_rs_1_10;
output 	io_w_dmem_dat_data_10;
output 	mem_rs_1_11;
output 	io_w_dmem_dat_data_11;
output 	mem_rs_1_12;
output 	io_w_dmem_dat_data_12;
output 	mem_rs_1_13;
output 	io_w_dmem_dat_data_13;
output 	mem_rs_1_14;
output 	io_w_dmem_dat_data_14;
output 	mem_rs_1_15;
output 	io_w_dmem_dat_data_15;
output 	mem_rs_1_16;
input 	data_out_17;
output 	mem_rs_1_17;
output 	mem_rs_1_18;
output 	mem_rs_1_19;
output 	mem_rs_1_20;
output 	mem_rs_1_21;
output 	mem_rs_1_22;
output 	mem_rs_1_23;
input 	data_out_27;
input 	av_readdata_pre_28;
input 	av_readdata_pre_29;
input 	av_readdata_pre_30;
input 	av_readdata_pre_31;
input 	av_readdata_pre_8;
input 	av_readdata_pre_9;
input 	av_readdata_pre_10;
input 	av_readdata_pre_11;
input 	av_readdata_pre_12;
input 	av_readdata_pre_13;
input 	av_readdata_pre_14;
input 	av_readdata_pre_15;
input 	av_readdata_pre_16;
input 	av_readdata_pre_17;
input 	av_readdata_pre_18;
input 	av_readdata_pre_19;
input 	av_readdata_pre_4;
input 	av_readdata_pre_2;
input 	av_readdata_pre_3;
input 	av_readdata_pre_5;
input 	av_readdata_pre_6;
input 	av_readdata_pre_7;
input 	av_readdata_pre_20;
input 	av_readdata_pre_21;
input 	av_readdata_pre_22;
input 	av_readdata_pre_23;
input 	av_readdata_pre_24;
input 	av_readdata_pre_25;
input 	av_readdata_pre_26;
input 	av_readdata_pre_27;
output 	mem_ctrl_mem_wr00;
output 	w_req;
output 	mem_ctrl_mem_wr01;
output 	io_imem_add_addr_2;
output 	io_imem_add_addr_3;
output 	io_imem_add_addr_4;
output 	io_imem_add_addr_5;
output 	io_imem_add_addr_6;
output 	io_imem_add_addr_7;
output 	io_imem_add_addr_8;
output 	io_imem_add_addr_9;
output 	io_imem_add_addr_10;
output 	io_imem_add_addr_11;
output 	io_imem_add_addr_12;
output 	io_imem_add_addr_13;
output 	io_imem_add_addr_14;
input 	read_latency_shift_reg_01;
output 	_GEN_73_0;
output 	io_w_dmem_dat_data_24;
output 	io_w_dmem_dat_data_25;
output 	io_w_dmem_dat_data_26;
output 	io_w_dmem_dat_data_27;
output 	io_w_dmem_dat_data_28;
output 	io_w_dmem_dat_data_29;
output 	io_w_dmem_dat_data_30;
output 	io_w_dmem_dat_data_31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



kyogenrv_fpga_KyogenRVCpu krv(
	.q_a_16(q_a_16),
	.q_a_15(q_a_15),
	.q_a_18(q_a_18),
	.q_a_17(q_a_17),
	.q_a_19(q_a_19),
	.q_a_21(q_a_21),
	.q_a_20(q_a_20),
	.q_a_23(q_a_23),
	.q_a_22(q_a_22),
	.q_a_24(q_a_24),
	.q_a_14(q_a_14),
	.q_a_13(q_a_13),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.q_a_12(q_a_12),
	.q_a_10(q_a_10),
	.q_a_11(q_a_11),
	.q_a_25(q_a_25),
	.q_a_30(q_a_30),
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_3(q_a_3),
	.q_a_2(q_a_2),
	.q_a_4(q_a_4),
	.q_a_26(q_a_26),
	.q_a_27(q_a_27),
	.q_a_31(q_a_31),
	.q_a_28(q_a_28),
	.q_a_29(q_a_29),
	.id_npc_0(id_npc_0),
	.id_npc_1(id_npc_1),
	.id_pc_2(id_pc_2),
	.id_pc_3(id_pc_3),
	.id_pc_4(id_pc_4),
	.id_pc_5(id_pc_5),
	.id_pc_6(id_pc_6),
	.id_pc_7(id_pc_7),
	.id_pc_8(id_pc_8),
	.id_pc_9(id_pc_9),
	.id_pc_10(id_pc_10),
	.id_pc_11(id_pc_11),
	.id_pc_12(id_pc_12),
	.id_pc_13(id_pc_13),
	.id_pc_14(id_pc_14),
	.id_pc_15(id_pc_15),
	.id_pc_16(id_pc_16),
	.id_pc_17(id_pc_17),
	.id_pc_18(id_pc_18),
	.id_pc_19(id_pc_19),
	.id_pc_20(id_pc_20),
	.id_pc_21(id_pc_21),
	.id_pc_22(id_pc_22),
	.id_pc_23(id_pc_23),
	.id_pc_24(id_pc_24),
	.id_pc_25(id_pc_25),
	.id_pc_26(id_pc_26),
	.id_pc_27(id_pc_27),
	.id_pc_28(id_pc_28),
	.id_pc_29(id_pc_29),
	.id_pc_30(id_pc_30),
	.id_pc_31(id_pc_31),
	.mem_alu_out_1(mem_alu_out_1),
	.av_readdata_pre_1(av_readdata_pre_1),
	.mem_alu_out_0(mem_alu_out_0),
	.av_readdata_pre_0(av_readdata_pre_0),
	.waitrequest_reset_override(waitrequest_reset_override),
	.wait_latency_counter_0(wait_latency_counter_0),
	.mem_ctrl_mem_wr10(mem_ctrl_mem_wr10),
	.wait_latency_counter_1(wait_latency_counter_1),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.mem_rs_1_0(mem_rs_1_0),
	.Equal68(Equal68),
	.Equal73(Equal73),
	.io_w_dmem_dat_data_0(io_w_dmem_dat_data_0),
	.mem_alu_out_2(mem_alu_out_2),
	.mem_alu_out_3(mem_alu_out_3),
	.mem_rs_1_1(mem_rs_1_1),
	.io_w_dmem_dat_data_1(io_w_dmem_dat_data_1),
	.mem_rs_1_2(mem_rs_1_2),
	.io_w_dmem_dat_data_2(io_w_dmem_dat_data_2),
	.mem_rs_1_3(mem_rs_1_3),
	.io_w_dmem_dat_data_3(io_w_dmem_dat_data_3),
	.mem_rs_1_4(mem_rs_1_4),
	.io_w_dmem_dat_data_4(io_w_dmem_dat_data_4),
	.mem_rs_1_5(mem_rs_1_5),
	.io_w_dmem_dat_data_5(io_w_dmem_dat_data_5),
	.mem_rs_1_6(mem_rs_1_6),
	.io_w_dmem_dat_data_6(io_w_dmem_dat_data_6),
	.mem_rs_1_7(mem_rs_1_7),
	.io_w_dmem_dat_data_7(io_w_dmem_dat_data_7),
	.mem_rs_1_8(mem_rs_1_8),
	.data_out_12(data_out_12),
	.io_w_dmem_dat_data_8(io_w_dmem_dat_data_8),
	.mem_rs_1_9(mem_rs_1_9),
	.io_w_dmem_dat_data_9(io_w_dmem_dat_data_9),
	.mem_rs_1_10(mem_rs_1_10),
	.io_w_dmem_dat_data_10(io_w_dmem_dat_data_10),
	.mem_rs_1_11(mem_rs_1_11),
	.io_w_dmem_dat_data_11(io_w_dmem_dat_data_11),
	.mem_rs_1_12(mem_rs_1_12),
	.io_w_dmem_dat_data_12(io_w_dmem_dat_data_12),
	.mem_rs_1_13(mem_rs_1_13),
	.io_w_dmem_dat_data_13(io_w_dmem_dat_data_13),
	.mem_rs_1_14(mem_rs_1_14),
	.io_w_dmem_dat_data_14(io_w_dmem_dat_data_14),
	.mem_rs_1_15(mem_rs_1_15),
	.io_w_dmem_dat_data_15(io_w_dmem_dat_data_15),
	.mem_rs_1_16(mem_rs_1_16),
	.data_out_17(data_out_17),
	.mem_rs_1_17(mem_rs_1_17),
	.mem_rs_1_18(mem_rs_1_18),
	.mem_rs_1_19(mem_rs_1_19),
	.mem_rs_1_20(mem_rs_1_20),
	.mem_rs_1_21(mem_rs_1_21),
	.mem_rs_1_22(mem_rs_1_22),
	.mem_rs_1_23(mem_rs_1_23),
	.data_out_27(data_out_27),
	.av_readdata_pre_28(av_readdata_pre_28),
	.av_readdata_pre_29(av_readdata_pre_29),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata_pre_31(av_readdata_pre_31),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_16(av_readdata_pre_16),
	.av_readdata_pre_17(av_readdata_pre_17),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_19(av_readdata_pre_19),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_2(av_readdata_pre_2),
	.av_readdata_pre_3(av_readdata_pre_3),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_6(av_readdata_pre_6),
	.av_readdata_pre_7(av_readdata_pre_7),
	.av_readdata_pre_20(av_readdata_pre_20),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_22(av_readdata_pre_22),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_24(av_readdata_pre_24),
	.av_readdata_pre_25(av_readdata_pre_25),
	.av_readdata_pre_26(av_readdata_pre_26),
	.av_readdata_pre_27(av_readdata_pre_27),
	.mem_ctrl_mem_wr00(mem_ctrl_mem_wr00),
	.w_req1(w_req),
	.mem_ctrl_mem_wr01(mem_ctrl_mem_wr01),
	.io_imem_add_addr_2(io_imem_add_addr_2),
	.io_imem_add_addr_3(io_imem_add_addr_3),
	.io_imem_add_addr_4(io_imem_add_addr_4),
	.io_imem_add_addr_5(io_imem_add_addr_5),
	.io_imem_add_addr_6(io_imem_add_addr_6),
	.io_imem_add_addr_7(io_imem_add_addr_7),
	.io_imem_add_addr_8(io_imem_add_addr_8),
	.io_imem_add_addr_9(io_imem_add_addr_9),
	.io_imem_add_addr_10(io_imem_add_addr_10),
	.io_imem_add_addr_11(io_imem_add_addr_11),
	.io_imem_add_addr_12(io_imem_add_addr_12),
	.io_imem_add_addr_13(io_imem_add_addr_13),
	.io_imem_add_addr_14(io_imem_add_addr_14),
	.read_latency_shift_reg_01(read_latency_shift_reg_01),
	._GEN_73_0(_GEN_73_0),
	.io_w_dmem_dat_data_24(io_w_dmem_dat_data_24),
	.io_w_dmem_dat_data_25(io_w_dmem_dat_data_25),
	.io_w_dmem_dat_data_26(io_w_dmem_dat_data_26),
	.io_w_dmem_dat_data_27(io_w_dmem_dat_data_27),
	.io_w_dmem_dat_data_28(io_w_dmem_dat_data_28),
	.io_w_dmem_dat_data_29(io_w_dmem_dat_data_29),
	.io_w_dmem_dat_data_30(io_w_dmem_dat_data_30),
	.io_w_dmem_dat_data_31(io_w_dmem_dat_data_31),
	.clk_clk(clk_clk));

endmodule

module kyogenrv_fpga_KyogenRVCpu (
	q_a_16,
	q_a_15,
	q_a_18,
	q_a_17,
	q_a_19,
	q_a_21,
	q_a_20,
	q_a_23,
	q_a_22,
	q_a_24,
	q_a_14,
	q_a_13,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	q_a_12,
	q_a_10,
	q_a_11,
	q_a_25,
	q_a_30,
	q_a_0,
	q_a_1,
	q_a_3,
	q_a_2,
	q_a_4,
	q_a_26,
	q_a_27,
	q_a_31,
	q_a_28,
	q_a_29,
	id_npc_0,
	id_npc_1,
	id_pc_2,
	id_pc_3,
	id_pc_4,
	id_pc_5,
	id_pc_6,
	id_pc_7,
	id_pc_8,
	id_pc_9,
	id_pc_10,
	id_pc_11,
	id_pc_12,
	id_pc_13,
	id_pc_14,
	id_pc_15,
	id_pc_16,
	id_pc_17,
	id_pc_18,
	id_pc_19,
	id_pc_20,
	id_pc_21,
	id_pc_22,
	id_pc_23,
	id_pc_24,
	id_pc_25,
	id_pc_26,
	id_pc_27,
	id_pc_28,
	id_pc_29,
	id_pc_30,
	id_pc_31,
	mem_alu_out_1,
	av_readdata_pre_1,
	mem_alu_out_0,
	av_readdata_pre_0,
	waitrequest_reset_override,
	wait_latency_counter_0,
	mem_ctrl_mem_wr10,
	wait_latency_counter_1,
	read_latency_shift_reg_0,
	altera_reset_synchronizer_int_chain_out,
	mem_rs_1_0,
	Equal68,
	Equal73,
	io_w_dmem_dat_data_0,
	mem_alu_out_2,
	mem_alu_out_3,
	mem_rs_1_1,
	io_w_dmem_dat_data_1,
	mem_rs_1_2,
	io_w_dmem_dat_data_2,
	mem_rs_1_3,
	io_w_dmem_dat_data_3,
	mem_rs_1_4,
	io_w_dmem_dat_data_4,
	mem_rs_1_5,
	io_w_dmem_dat_data_5,
	mem_rs_1_6,
	io_w_dmem_dat_data_6,
	mem_rs_1_7,
	io_w_dmem_dat_data_7,
	mem_rs_1_8,
	data_out_12,
	io_w_dmem_dat_data_8,
	mem_rs_1_9,
	io_w_dmem_dat_data_9,
	mem_rs_1_10,
	io_w_dmem_dat_data_10,
	mem_rs_1_11,
	io_w_dmem_dat_data_11,
	mem_rs_1_12,
	io_w_dmem_dat_data_12,
	mem_rs_1_13,
	io_w_dmem_dat_data_13,
	mem_rs_1_14,
	io_w_dmem_dat_data_14,
	mem_rs_1_15,
	io_w_dmem_dat_data_15,
	mem_rs_1_16,
	data_out_17,
	mem_rs_1_17,
	mem_rs_1_18,
	mem_rs_1_19,
	mem_rs_1_20,
	mem_rs_1_21,
	mem_rs_1_22,
	mem_rs_1_23,
	data_out_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_30,
	av_readdata_pre_31,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata_pre_18,
	av_readdata_pre_19,
	av_readdata_pre_4,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_20,
	av_readdata_pre_21,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_27,
	mem_ctrl_mem_wr00,
	w_req1,
	mem_ctrl_mem_wr01,
	io_imem_add_addr_2,
	io_imem_add_addr_3,
	io_imem_add_addr_4,
	io_imem_add_addr_5,
	io_imem_add_addr_6,
	io_imem_add_addr_7,
	io_imem_add_addr_8,
	io_imem_add_addr_9,
	io_imem_add_addr_10,
	io_imem_add_addr_11,
	io_imem_add_addr_12,
	io_imem_add_addr_13,
	io_imem_add_addr_14,
	read_latency_shift_reg_01,
	_GEN_73_0,
	io_w_dmem_dat_data_24,
	io_w_dmem_dat_data_25,
	io_w_dmem_dat_data_26,
	io_w_dmem_dat_data_27,
	io_w_dmem_dat_data_28,
	io_w_dmem_dat_data_29,
	io_w_dmem_dat_data_30,
	io_w_dmem_dat_data_31,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	q_a_16;
input 	q_a_15;
input 	q_a_18;
input 	q_a_17;
input 	q_a_19;
input 	q_a_21;
input 	q_a_20;
input 	q_a_23;
input 	q_a_22;
input 	q_a_24;
input 	q_a_14;
input 	q_a_13;
input 	q_a_5;
input 	q_a_6;
input 	q_a_7;
input 	q_a_8;
input 	q_a_9;
input 	q_a_12;
input 	q_a_10;
input 	q_a_11;
input 	q_a_25;
input 	q_a_30;
input 	q_a_0;
input 	q_a_1;
input 	q_a_3;
input 	q_a_2;
input 	q_a_4;
input 	q_a_26;
input 	q_a_27;
input 	q_a_31;
input 	q_a_28;
input 	q_a_29;
output 	id_npc_0;
output 	id_npc_1;
output 	id_pc_2;
output 	id_pc_3;
output 	id_pc_4;
output 	id_pc_5;
output 	id_pc_6;
output 	id_pc_7;
output 	id_pc_8;
output 	id_pc_9;
output 	id_pc_10;
output 	id_pc_11;
output 	id_pc_12;
output 	id_pc_13;
output 	id_pc_14;
output 	id_pc_15;
output 	id_pc_16;
output 	id_pc_17;
output 	id_pc_18;
output 	id_pc_19;
output 	id_pc_20;
output 	id_pc_21;
output 	id_pc_22;
output 	id_pc_23;
output 	id_pc_24;
output 	id_pc_25;
output 	id_pc_26;
output 	id_pc_27;
output 	id_pc_28;
output 	id_pc_29;
output 	id_pc_30;
output 	id_pc_31;
output 	mem_alu_out_1;
input 	av_readdata_pre_1;
output 	mem_alu_out_0;
input 	av_readdata_pre_0;
input 	waitrequest_reset_override;
input 	wait_latency_counter_0;
output 	mem_ctrl_mem_wr10;
input 	wait_latency_counter_1;
input 	read_latency_shift_reg_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	mem_rs_1_0;
output 	Equal68;
output 	Equal73;
output 	io_w_dmem_dat_data_0;
output 	mem_alu_out_2;
output 	mem_alu_out_3;
output 	mem_rs_1_1;
output 	io_w_dmem_dat_data_1;
output 	mem_rs_1_2;
output 	io_w_dmem_dat_data_2;
output 	mem_rs_1_3;
output 	io_w_dmem_dat_data_3;
output 	mem_rs_1_4;
output 	io_w_dmem_dat_data_4;
output 	mem_rs_1_5;
output 	io_w_dmem_dat_data_5;
output 	mem_rs_1_6;
output 	io_w_dmem_dat_data_6;
output 	mem_rs_1_7;
output 	io_w_dmem_dat_data_7;
output 	mem_rs_1_8;
input 	data_out_12;
output 	io_w_dmem_dat_data_8;
output 	mem_rs_1_9;
output 	io_w_dmem_dat_data_9;
output 	mem_rs_1_10;
output 	io_w_dmem_dat_data_10;
output 	mem_rs_1_11;
output 	io_w_dmem_dat_data_11;
output 	mem_rs_1_12;
output 	io_w_dmem_dat_data_12;
output 	mem_rs_1_13;
output 	io_w_dmem_dat_data_13;
output 	mem_rs_1_14;
output 	io_w_dmem_dat_data_14;
output 	mem_rs_1_15;
output 	io_w_dmem_dat_data_15;
output 	mem_rs_1_16;
input 	data_out_17;
output 	mem_rs_1_17;
output 	mem_rs_1_18;
output 	mem_rs_1_19;
output 	mem_rs_1_20;
output 	mem_rs_1_21;
output 	mem_rs_1_22;
output 	mem_rs_1_23;
input 	data_out_27;
input 	av_readdata_pre_28;
input 	av_readdata_pre_29;
input 	av_readdata_pre_30;
input 	av_readdata_pre_31;
input 	av_readdata_pre_8;
input 	av_readdata_pre_9;
input 	av_readdata_pre_10;
input 	av_readdata_pre_11;
input 	av_readdata_pre_12;
input 	av_readdata_pre_13;
input 	av_readdata_pre_14;
input 	av_readdata_pre_15;
input 	av_readdata_pre_16;
input 	av_readdata_pre_17;
input 	av_readdata_pre_18;
input 	av_readdata_pre_19;
input 	av_readdata_pre_4;
input 	av_readdata_pre_2;
input 	av_readdata_pre_3;
input 	av_readdata_pre_5;
input 	av_readdata_pre_6;
input 	av_readdata_pre_7;
input 	av_readdata_pre_20;
input 	av_readdata_pre_21;
input 	av_readdata_pre_22;
input 	av_readdata_pre_23;
input 	av_readdata_pre_24;
input 	av_readdata_pre_25;
input 	av_readdata_pre_26;
input 	av_readdata_pre_27;
output 	mem_ctrl_mem_wr00;
output 	w_req1;
output 	mem_ctrl_mem_wr01;
output 	io_imem_add_addr_2;
output 	io_imem_add_addr_3;
output 	io_imem_add_addr_4;
output 	io_imem_add_addr_5;
output 	io_imem_add_addr_6;
output 	io_imem_add_addr_7;
output 	io_imem_add_addr_8;
output 	io_imem_add_addr_9;
output 	io_imem_add_addr_10;
output 	io_imem_add_addr_11;
output 	io_imem_add_addr_12;
output 	io_imem_add_addr_13;
output 	io_imem_add_addr_14;
input 	read_latency_shift_reg_01;
output 	_GEN_73_0;
output 	io_w_dmem_dat_data_24;
output 	io_w_dmem_dat_data_25;
output 	io_w_dmem_dat_data_26;
output 	io_w_dmem_dat_data_27;
output 	io_w_dmem_dat_data_28;
output 	io_w_dmem_dat_data_29;
output 	io_w_dmem_dat_data_30;
output 	io_w_dmem_dat_data_31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ex_j_check~q ;
wire \_T_3549~q ;
wire \alu|_T_3[0]~0_combout ;
wire \alu|_T_3[1]~2_combout ;
wire \alu|_T_3[2]~4_combout ;
wire \alu|_T_3[3]~6_combout ;
wire \alu|_T_3[4]~8_combout ;
wire \alu|_T_3[5]~10_combout ;
wire \alu|_T_3[6]~12_combout ;
wire \alu|_T_3[7]~14_combout ;
wire \alu|_T_3[8]~16_combout ;
wire \alu|_T_3[9]~18_combout ;
wire \alu|_T_3[10]~20_combout ;
wire \alu|_T_3[11]~22_combout ;
wire \alu|_T_3[12]~24_combout ;
wire \alu|_T_3[13]~26_combout ;
wire \alu|_T_3[14]~28_combout ;
wire \alu|_T_3[15]~30_combout ;
wire \alu|_T_3[16]~32_combout ;
wire \alu|_T_3[17]~34_combout ;
wire \alu|_T_3[18]~36_combout ;
wire \alu|_T_3[19]~38_combout ;
wire \alu|_T_3[20]~40_combout ;
wire \alu|_T_3[21]~42_combout ;
wire \alu|_T_3[22]~44_combout ;
wire \alu|_T_3[23]~46_combout ;
wire \alu|_T_3[24]~48_combout ;
wire \alu|_T_3[25]~50_combout ;
wire \alu|_T_3[26]~52_combout ;
wire \alu|_T_3[27]~54_combout ;
wire \alu|_T_3[28]~56_combout ;
wire \alu|_T_3[29]~58_combout ;
wire \alu|_T_3[30]~60_combout ;
wire \alu|_T_3[31]~62_combout ;
wire \csr|mepc[2]~q ;
wire \csr|mepc[3]~q ;
wire \csr|mepc[4]~q ;
wire \csr|mepc[5]~q ;
wire \csr|mepc[6]~q ;
wire \csr|mepc[7]~q ;
wire \csr|mepc[8]~q ;
wire \csr|mepc[9]~q ;
wire \csr|mepc[10]~q ;
wire \csr|mepc[11]~q ;
wire \csr|mepc[12]~q ;
wire \csr|mepc[13]~q ;
wire \csr|mepc[14]~q ;
wire \csr|mepc[15]~q ;
wire \csr|mepc[16]~q ;
wire \csr|mepc[17]~q ;
wire \csr|mepc[18]~q ;
wire \csr|mepc[19]~q ;
wire \csr|mepc[20]~q ;
wire \csr|mepc[21]~q ;
wire \csr|mepc[22]~q ;
wire \csr|mepc[23]~q ;
wire \csr|mepc[24]~q ;
wire \csr|mepc[25]~q ;
wire \csr|mepc[26]~q ;
wire \csr|mepc[27]~q ;
wire \csr|mepc[28]~q ;
wire \csr|mepc[29]~q ;
wire \csr|mepc[30]~q ;
wire \csr|mepc[31]~q ;
wire \ex_b_check~q ;
wire \Equal56~0_combout ;
wire \Equal56~1_combout ;
wire \Equal56~2_combout ;
wire \Equal56~3_combout ;
wire \Equal56~4_combout ;
wire \Equal56~5_combout ;
wire \Equal56~6_combout ;
wire \Equal56~7_combout ;
wire \Equal56~8_combout ;
wire \Equal56~9_combout ;
wire \Equal56~10_combout ;
wire \ex_ctrl_legal~q ;
wire \csr_io_alu_op1[0]~4_combout ;
wire \csr|io_expt~0_combout ;
wire \_T_3557~0_combout ;
wire \_T_3557~1_combout ;
wire \_T_3557~2_combout ;
wire \_T_3557~3_combout ;
wire \_T_3557~4_combout ;
wire \_T_3557~5_combout ;
wire \_T_3557~6_combout ;
wire \csr|mcause[0]~6_combout ;
wire \ex_csr_cmd[2]~q ;
wire \ex_csr_cmd[0]~q ;
wire \ex_csr_cmd[1]~q ;
wire \csr|isEcall~0_combout ;
wire \csr|mepc[0]~q ;
wire \csr|io_expt~combout ;
wire \csr|mtvec[0]~q ;
wire \alu|_T_123[31]~combout ;
wire \alu|_T_123[11]~combout ;
wire \alu|_T_123[15]~combout ;
wire \alu|_T_123[19]~combout ;
wire \alu|_T_123[2]~combout ;
wire \alu|_T_123[7]~combout ;
wire \alu_io_op1[23]~60_combout ;
wire \alu_io_op1[27]~61_combout ;
wire \alu|LessThan0~0_combout ;
wire \alu|_T_125~20_combout ;
wire \ex_ctrl_legal~2_combout ;
wire \_GEN_32~0_combout ;
wire \_GEN_32~1_combout ;
wire \alu_io_op1[31]~62_combout ;
wire \csr_io_alu_op1[0]~5_combout ;
wire \alu_io_op1[30]~63_combout ;
wire \csr_io_alu_op1[1]~6_combout ;
wire \alu|ShiftRight0~38_combout ;
wire \alu_io_op1[8]~64_combout ;
wire \alu_io_op1[7]~65_combout ;
wire \alu_io_op1[24]~66_combout ;
wire \alu_io_op1[4]~67_combout ;
wire \alu_io_op1[3]~68_combout ;
wire \alu_io_op1[28]~69_combout ;
wire \alu_io_op1[6]~70_combout ;
wire \alu_io_op1[25]~71_combout ;
wire \alu_io_op1[5]~72_combout ;
wire \alu_io_op1[26]~73_combout ;
wire \alu_io_op1[2]~74_combout ;
wire \alu_io_op1[29]~75_combout ;
wire \alu_io_op1[12]~76_combout ;
wire \alu_io_op1[19]~77_combout ;
wire \alu_io_op1[11]~78_combout ;
wire \alu_io_op1[20]~79_combout ;
wire \alu_io_op1[10]~80_combout ;
wire \alu_io_op1[21]~81_combout ;
wire \alu_io_op1[9]~82_combout ;
wire \alu_io_op1[22]~83_combout ;
wire \alu_io_op1[16]~84_combout ;
wire \alu_io_op1[15]~85_combout ;
wire \alu_io_op1[14]~86_combout ;
wire \alu_io_op1[17]~87_combout ;
wire \alu_io_op1[13]~88_combout ;
wire \alu_io_op1[18]~89_combout ;
wire \alu|ShiftRight0~94_combout ;
wire \csr|mepc[1]~q ;
wire \csr|mtvec[1]~q ;
wire \csr|io_out[1]~16_combout ;
wire \csr|io_out[0]~24_combout ;
wire \alu|ShiftRight0~126_combout ;
wire \alu|ShiftRight0~128_combout ;
wire \alu|io_out[0]~1_combout ;
wire \wb_dmem_read_ack~q ;
wire \_GEN_9~combout ;
wire \ex_ctrl_csr_cmd~15_combout ;
wire \Equal47~0_combout ;
wire \ex_csr_cmd~6_combout ;
wire \ex_csr_cmd~7_combout ;
wire \ex_csr_cmd~8_combout ;
wire \ex_csr_cmd~9_combout ;
wire \csr|mtvec[2]~q ;
wire \csr|mtvec[3]~q ;
wire \csr|mtvec[4]~q ;
wire \csr|mtvec[5]~q ;
wire \csr|mtvec[6]~q ;
wire \csr|mtvec[7]~q ;
wire \csr|mtvec[8]~q ;
wire \csr|mtvec[9]~q ;
wire \csr|mtvec[10]~q ;
wire \csr|mtvec[11]~q ;
wire \csr|mtvec[12]~q ;
wire \csr|mtvec[13]~q ;
wire \csr|mtvec[14]~q ;
wire \csr|mtvec[15]~q ;
wire \csr|mtvec[16]~q ;
wire \csr|mtvec[17]~q ;
wire \csr|mtvec[18]~q ;
wire \csr|mtvec[19]~q ;
wire \csr|mtvec[20]~q ;
wire \csr|mtvec[21]~q ;
wire \csr|mtvec[22]~q ;
wire \csr|mtvec[23]~q ;
wire \csr|mtvec[24]~q ;
wire \csr|mtvec[25]~q ;
wire \csr|mtvec[26]~q ;
wire \csr|mtvec[27]~q ;
wire \csr|mtvec[28]~q ;
wire \csr|mtvec[29]~q ;
wire \csr|mtvec[30]~q ;
wire \csr|mtvec[31]~q ;
wire \alu|ShiftRight0~130_combout ;
wire \alu|ShiftRight0~150_combout ;
wire \alu|ShiftRight0~152_combout ;
wire \alu|ShiftRight0~167_combout ;
wire \io_sw_r_ex_imm[0]~9_combout ;
wire \csr_io_in[0]~1_combout ;
wire \csr_io_in[0]~2_combout ;
wire \csr_io_in[0]~3_combout ;
wire \csr_io_in[0]~4_combout ;
wire \csr_io_in[0]~5_combout ;
wire \csr_io_in[0]~6_combout ;
wire \csr|io_out[28]~31_combout ;
wire \csr|io_out[29]~36_combout ;
wire \csr|io_out[29]~37_combout ;
wire \csr|io_out[30]~45_combout ;
wire \csr|io_out[31]~52_combout ;
wire \alu|ShiftRight0~173_combout ;
wire \alu|ShiftRight0~175_combout ;
wire \csr|io_out[8]~59_combout ;
wire \alu|ShiftRight0~180_combout ;
wire \alu|ShiftRight0~183_combout ;
wire \csr|io_out[9]~66_combout ;
wire \alu|ShiftRight0~188_combout ;
wire \alu|ShiftRight0~190_combout ;
wire \csr|io_out[10]~72_combout ;
wire \alu|ShiftRight0~195_combout ;
wire \alu|ShiftRight0~197_combout ;
wire \csr|io_out[11]~79_combout ;
wire \alu|ShiftRight0~198_combout ;
wire \alu|ShiftRight0~203_combout ;
wire \csr|io_out[12]~86_combout ;
wire \alu|_T_123[13]~combout ;
wire \alu|ShiftRight0~209_combout ;
wire \csr|io_out[13]~93_combout ;
wire \alu|ShiftRight0~216_combout ;
wire \csr|io_out[14]~100_combout ;
wire \alu|ShiftRight0~217_combout ;
wire \alu|ShiftRight0~222_combout ;
wire \csr|io_out[15]~107_combout ;
wire \csr|io_out[16]~114_combout ;
wire \csr|io_out[17]~121_combout ;
wire \csr|io_out[18]~128_combout ;
wire \alu|_T_139[18]~combout ;
wire \csr|io_out[19]~135_combout ;
wire \csr|io_out[4]~142_combout ;
wire \alu|ShiftRight0~228_combout ;
wire \csr|io_out[2]~150_combout ;
wire \csr|io_out[3]~159_combout ;
wire \alu|ShiftRight0~233_combout ;
wire \csr|io_out[5]~166_combout ;
wire \alu|ShiftRight0~236_combout ;
wire \csr|io_out[6]~173_combout ;
wire \alu|ShiftRight0~240_combout ;
wire \csr|io_out[7]~181_combout ;
wire \csr|io_out[20]~188_combout ;
wire \csr|io_out[21]~193_combout ;
wire \csr|io_out[21]~194_combout ;
wire \csr|io_out[22]~202_combout ;
wire \csr|io_out[23]~209_combout ;
wire \csr|io_out[24]~216_combout ;
wire \csr|io_out[25]~221_combout ;
wire \csr|io_out[25]~222_combout ;
wire \csr|io_out[26]~230_combout ;
wire \csr|io_out[27]~235_combout ;
wire \csr|io_out[27]~236_combout ;
wire \csr_io_in[1]~7_combout ;
wire \csr_io_in[1]~8_combout ;
wire \csr_io_in[1]~9_combout ;
wire \csr_io_in[1]~10_combout ;
wire \ex_inst[0]~q ;
wire \ex_inst[1]~q ;
wire \ex_inst[4]~q ;
wire \ex_inst[2]~q ;
wire \ex_inst[3]~q ;
wire \ex_inst[5]~q ;
wire \ex_inst[6]~q ;
wire \wb_dmem_read_ack~0_combout ;
wire \csr_io_in[2]~11_combout ;
wire \csr_io_in[2]~12_combout ;
wire \csr_io_in[2]~13_combout ;
wire \csr_io_in[2]~14_combout ;
wire \csr_io_in[3]~15_combout ;
wire \csr_io_in[3]~16_combout ;
wire \csr_io_in[3]~17_combout ;
wire \csr_io_in[3]~18_combout ;
wire \csr_io_in[4]~19_combout ;
wire \csr_io_in[4]~20_combout ;
wire \csr_io_in[4]~21_combout ;
wire \csr_io_in[4]~22_combout ;
wire \csr_io_in[5]~23_combout ;
wire \csr_io_in[5]~24_combout ;
wire \csr_io_in[5]~25_combout ;
wire \csr_io_in[6]~26_combout ;
wire \csr_io_in[6]~27_combout ;
wire \csr_io_in[6]~28_combout ;
wire \csr_io_in[7]~29_combout ;
wire \csr_io_in[7]~30_combout ;
wire \csr_io_in[7]~31_combout ;
wire \csr_io_in[8]~32_combout ;
wire \csr_io_in[8]~33_combout ;
wire \csr_io_in[8]~34_combout ;
wire \csr_io_in[9]~35_combout ;
wire \csr_io_in[9]~36_combout ;
wire \csr_io_in[9]~37_combout ;
wire \csr_io_in[10]~38_combout ;
wire \csr_io_in[10]~39_combout ;
wire \csr_io_in[10]~40_combout ;
wire \csr_io_in[11]~41_combout ;
wire \csr_io_in[11]~42_combout ;
wire \csr_io_in[11]~43_combout ;
wire \csr_io_in[12]~44_combout ;
wire \csr_io_in[12]~45_combout ;
wire \csr_io_in[12]~46_combout ;
wire \csr_io_in[13]~47_combout ;
wire \csr_io_in[13]~48_combout ;
wire \csr_io_in[13]~49_combout ;
wire \csr_io_in[14]~50_combout ;
wire \csr_io_in[14]~51_combout ;
wire \csr_io_in[14]~52_combout ;
wire \csr_io_in[15]~53_combout ;
wire \csr_io_in[15]~54_combout ;
wire \csr_io_in[15]~55_combout ;
wire \csr_io_in[16]~56_combout ;
wire \csr_io_in[16]~57_combout ;
wire \csr_io_in[16]~58_combout ;
wire \csr_io_in[17]~59_combout ;
wire \csr_io_in[17]~60_combout ;
wire \csr_io_in[17]~61_combout ;
wire \csr_io_in[18]~62_combout ;
wire \csr_io_in[18]~63_combout ;
wire \csr_io_in[18]~64_combout ;
wire \csr_io_in[19]~65_combout ;
wire \csr_io_in[19]~66_combout ;
wire \csr_io_in[19]~67_combout ;
wire \csr_io_in[20]~68_combout ;
wire \csr_io_in[20]~69_combout ;
wire \csr_io_in[20]~70_combout ;
wire \csr_io_in[21]~71_combout ;
wire \csr_io_in[21]~72_combout ;
wire \csr_io_in[21]~73_combout ;
wire \csr_io_in[22]~74_combout ;
wire \csr_io_in[22]~75_combout ;
wire \csr_io_in[22]~76_combout ;
wire \csr_io_in[23]~77_combout ;
wire \csr_io_in[23]~78_combout ;
wire \csr_io_in[23]~79_combout ;
wire \csr_io_in[24]~80_combout ;
wire \csr_io_in[24]~81_combout ;
wire \csr_io_in[24]~82_combout ;
wire \csr_io_in[25]~83_combout ;
wire \csr_io_in[25]~84_combout ;
wire \csr_io_in[25]~85_combout ;
wire \csr_io_in[26]~86_combout ;
wire \csr_io_in[26]~87_combout ;
wire \csr_io_in[26]~88_combout ;
wire \csr_io_in[27]~89_combout ;
wire \csr_io_in[27]~90_combout ;
wire \csr_io_in[27]~91_combout ;
wire \csr_io_in[28]~92_combout ;
wire \csr_io_in[28]~93_combout ;
wire \csr_io_in[28]~94_combout ;
wire \csr_io_in[29]~95_combout ;
wire \csr_io_in[29]~96_combout ;
wire \csr_io_in[29]~97_combout ;
wire \csr_io_in[30]~98_combout ;
wire \csr_io_in[30]~99_combout ;
wire \csr_io_in[30]~100_combout ;
wire \csr_io_in[31]~101_combout ;
wire \csr_io_in[31]~102_combout ;
wire \csr_io_in[31]~103_combout ;
wire \csr_io_in[31]~104_combout ;
wire \ex_inst~13_combout ;
wire \ex_inst~14_combout ;
wire \ex_inst~15_combout ;
wire \ex_inst~16_combout ;
wire \ex_inst~17_combout ;
wire \ex_inst~18_combout ;
wire \ex_inst~19_combout ;
wire \alu|_T_123[23]~combout ;
wire \alu|_T_123[27]~combout ;
wire \ex_ctrl_legal~3_combout ;
wire \alu|_T_123[29]~combout ;
wire \alu|ShiftRight0~249_combout ;
wire \alu|ShiftRight0~250_combout ;
wire \alu|_T_123[17]~combout ;
wire \alu|ShiftRight0~251_combout ;
wire \alu|ShiftRight0~253_combout ;
wire \alu|ShiftRight0~254_combout ;
wire \alu|ShiftRight0~256_combout ;
wire \alu|_T_123[21]~combout ;
wire \alu|_T_123[25]~combout ;
wire \_GEN_33~2_combout ;
wire \_T_1778~combout ;
wire \id_inst~21_combout ;
wire \id_inst~0_combout ;
wire \id_pc[7]~0_combout ;
wire \id_inst[14]~q ;
wire \id_inst~33_combout ;
wire \id_inst[0]~q ;
wire \id_inst~34_combout ;
wire \id_inst[1]~q ;
wire \id_inst~35_combout ;
wire \id_inst[3]~q ;
wire \id_inst~36_combout ;
wire \id_inst[2]~q ;
wire \ex_ctrl_mem_wr~7_combout ;
wire \id_inst~23_combout ;
wire \id_inst[5]~q ;
wire \id_inst~24_combout ;
wire \id_inst[6]~q ;
wire \Equal7~0_combout ;
wire \id_inst~37_combout ;
wire \id_inst[4]~q ;
wire \Equal11~0_combout ;
wire \id_inst~28_combout ;
wire \id_inst[12]~q ;
wire \id_inst~22_combout ;
wire \id_inst[13]~q ;
wire \Equal14~0_combout ;
wire \Equal9~0_combout ;
wire \Equal8~1_combout ;
wire \Equal8~0_combout ;
wire \Equal10~0_combout ;
wire \Equal10~1_combout ;
wire \ex_ctrl_alu_func~4_combout ;
wire \id_ctrl_br_type[2]~11_combout ;
wire \Equal5~0_combout ;
wire \Equal8~2_combout ;
wire \_GEN_15~0_combout ;
wire \Equal53~0_combout ;
wire \Equal6~3_combout ;
wire \ex_ctrl_alu_op1~2_combout ;
wire \Equal5~1_combout ;
wire \ex_ctrl_imm_type~14_combout ;
wire \id_ctrl_br_type[0]~4_combout ;
wire \id_ctrl_br_type[2]~5_combout ;
wire \ex_ctrl_br_type~0_combout ;
wire \ex_ctrl_br_type[2]~q ;
wire \mem_ctrl_br_type~0_combout ;
wire \mem_ctrl_br_type[2]~q ;
wire \id_pc[7]~31_combout ;
wire \ex_ctrl_br_type~1_combout ;
wire \ex_ctrl_br_type[3]~q ;
wire \mem_ctrl_br_type~1_combout ;
wire \mem_ctrl_br_type[3]~q ;
wire \Equal2~0_combout ;
wire \id_inst~11_combout ;
wire \id_inst~12_combout ;
wire \id_inst[21]~q ;
wire \id_inst~3_combout ;
wire \id_inst~4_combout ;
wire \id_inst[15]~q ;
wire \id_inst~1_combout ;
wire \id_inst~2_combout ;
wire \id_inst[16]~q ;
wire \id_inst~7_combout ;
wire \id_inst~8_combout ;
wire \id_inst[17]~q ;
wire \id_inst~5_combout ;
wire \id_inst~6_combout ;
wire \id_inst[18]~q ;
wire \ex_rs_0[3]~0_combout ;
wire \id_inst~9_combout ;
wire \id_inst~10_combout ;
wire \id_inst[19]~q ;
wire \ex_rs_0[3]~1_combout ;
wire \id_inst~19_combout ;
wire \id_inst~20_combout ;
wire \id_inst[24]~q ;
wire \id_inst~17_combout ;
wire \id_inst~18_combout ;
wire \id_inst[22]~q ;
wire \id_inst~15_combout ;
wire \id_inst~16_combout ;
wire \id_inst[23]~q ;
wire \id_inst~25_combout ;
wire \id_inst[7]~q ;
wire \Equal48~0_combout ;
wire \id_inst~26_combout ;
wire \id_inst[8]~q ;
wire \id_inst~27_combout ;
wire \id_inst[9]~q ;
wire \Equal48~1_combout ;
wire \id_inst~29_combout ;
wire \id_inst[10]~q ;
wire \id_inst~30_combout ;
wire \id_inst[11]~q ;
wire \id_inst~31_combout ;
wire \id_inst[25]~q ;
wire \Equal48~2_combout ;
wire \id_inst~32_combout ;
wire \id_inst[30]~q ;
wire \Equal48~3_combout ;
wire \id_inst~38_combout ;
wire \id_inst[26]~q ;
wire \id_inst~39_combout ;
wire \id_inst[27]~q ;
wire \id_inst~40_combout ;
wire \id_inst[31]~q ;
wire \Equal49~0_combout ;
wire \id_inst~41_combout ;
wire \id_inst[28]~q ;
wire \id_inst~13_combout ;
wire \id_inst~14_combout ;
wire \id_inst[20]~q ;
wire \Equal49~1_combout ;
wire \Equal49~2_combout ;
wire \id_inst~42_combout ;
wire \id_inst[29]~q ;
wire \Equal49~3_combout ;
wire \Equal15~0_combout ;
wire \Equal17~0_combout ;
wire \Equal20~0_combout ;
wire \ex_ctrl_imm_type~11_combout ;
wire \Equal22~0_combout ;
wire \ex_ctrl_imm_type~12_combout ;
wire \Equal16~0_combout ;
wire \ex_ctrl_mask_type~1_combout ;
wire \Equal18~1_combout ;
wire \ex_ctrl_mask_type~2_combout ;
wire \Equal15~1_combout ;
wire \_T_3091~0_combout ;
wire \Equal6~2_combout ;
wire \ex_ctrl_alu_func~9_combout ;
wire \_T_2062[1]~0_combout ;
wire \id_ctrl_br_type[1]~6_combout ;
wire \id_ctrl_br_type[1]~12_combout ;
wire \id_ctrl_br_type[1]~10_combout ;
wire \ex_ctrl_br_type[1]~q ;
wire \mem_ctrl_br_type~3_combout ;
wire \mem_ctrl_br_type[1]~q ;
wire \inst_kill~1_combout ;
wire \Equal9~1_combout ;
wire \ex_ctrl_alu_func~10_combout ;
wire \Equal26~0_combout ;
wire \Equal13~0_combout ;
wire \Equal27~0_combout ;
wire \ex_ctrl_alu_func~34_combout ;
wire \Equal28~0_combout ;
wire \Equal28~1_combout ;
wire \Equal12~0_combout ;
wire \Equal29~0_combout ;
wire \Equal32~0_combout ;
wire \Equal39~0_combout ;
wire \Equal34~0_combout ;
wire \Equal37~0_combout ;
wire \ex_ctrl_alu_func~11_combout ;
wire \Equal18~0_combout ;
wire \Equal29~1_combout ;
wire \Equal31~0_combout ;
wire \Equal31~1_combout ;
wire \ex_ctrl_alu_op2~5_combout ;
wire \ex_ctrl_alu_func~12_combout ;
wire \ex_ctrl_alu_func~13_combout ;
wire \ex_ctrl_alu_func~14_combout ;
wire \ex_ctrl_alu_func~15_combout ;
wire \ex_ctrl_alu_func[0]~q ;
wire \_GEN_53~combout ;
wire \mem_alu_cmp_out~q ;
wire \inst_kill~0_combout ;
wire \mem_ctrl_mem_wr~7_combout ;
wire \id_ctrl_br_type[0]~7_combout ;
wire \id_ctrl_br_type[0]~8_combout ;
wire \id_ctrl_br_type[0]~9_combout ;
wire \ex_ctrl_br_type[0]~q ;
wire \mem_ctrl_br_type~2_combout ;
wire \mem_ctrl_br_type[0]~q ;
wire \Equal4~0_combout ;
wire \pc_cntr[0]~0_combout ;
wire \ex_inst~6_combout ;
wire \ex_inst[7]~q ;
wire \ex_inst~0_combout ;
wire \ex_inst[15]~q ;
wire \ex_ctrl_mask_type~0_combout ;
wire \ex_ctrl_alu_func~6_combout ;
wire \ex_ctrl_alu_func~7_combout ;
wire \_T_3083~0_combout ;
wire \ex_ctrl_alu_func~33_combout ;
wire \_GEN_15~1_combout ;
wire \_GEN_15~2_combout ;
wire \ex_ctrl_csr_cmd~9_combout ;
wire \Equal43~0_combout ;
wire \ex_ctrl_imm_type~13_combout ;
wire \ex_ctrl_imm_type~17_combout ;
wire \ex_ctrl_imm_type.101~q ;
wire \ex_csr_addr~0_combout ;
wire \ex_csr_addr[0]~q ;
wire \ex_ctrl_imm_type~18_combout ;
wire \ex_ctrl_imm_type~19_combout ;
wire \ex_csr_cmd~10_combout ;
wire \Equal32~1_combout ;
wire \Equal33~0_combout ;
wire \ex_ctrl_alu_func~8_combout ;
wire \Equal32~2_combout ;
wire \ex_ctrl_csr_cmd~10_combout ;
wire \ex_ctrl_csr_cmd~14_combout ;
wire \ex_ctrl_imm_type~20_combout ;
wire \ex_ctrl_imm_type.000~q ;
wire \io_sw_r_ex_imm[0]~2_combout ;
wire \ex_csr_cmd~5_combout ;
wire \ex_ctrl_mem_wr~8_combout ;
wire \ex_ctrl_mem_wr~9_combout ;
wire \ex_ctrl_mask_type~3_combout ;
wire \ex_ctrl_mem_wr~10_combout ;
wire \ex_ctrl_imm_type.001~q ;
wire \mem_imm~46_combout ;
wire \mem_imm[0]~q ;
wire \_T_3862[0]~0_combout ;
wire \pc_cntr[0]~1_combout ;
wire \pc_cntr~2_combout ;
wire \pc_cntr~3_combout ;
wire \pc_cntr[0]~4_combout ;
wire \pc_cntr[0]~q ;
wire \id_npc~0_combout ;
wire \ex_inst~5_combout ;
wire \ex_inst[8]~q ;
wire \ex_inst~1_combout ;
wire \ex_inst[16]~q ;
wire \ex_csr_addr~1_combout ;
wire \ex_csr_addr[1]~q ;
wire \io_sw_r_ex_imm[1]~0_combout ;
wire \ex_ctrl_alu_op1~3_combout ;
wire \ex_ctrl_imm_type~15_combout ;
wire \ex_ctrl_imm_type.010~q ;
wire \io_sw_r_ex_imm[1]~1_combout ;
wire \ex_ctrl_imm_type~16_combout ;
wire \ex_ctrl_imm_type.011~q ;
wire \mem_imm~16_combout ;
wire \mem_imm[1]~q ;
wire \_T_3862[1]~2_combout ;
wire \pc_cntr~5_combout ;
wire \pc_cntr~6_combout ;
wire \pc_cntr[1]~q ;
wire \id_npc~1_combout ;
wire \ex_pc~4_combout ;
wire \ex_pc[2]~q ;
wire \mem_pc~0_combout ;
wire \mem_pc[2]~q ;
wire \ex_inst~7_combout ;
wire \ex_inst[9]~q ;
wire \ex_inst~2_combout ;
wire \ex_inst[17]~q ;
wire \ex_csr_addr~2_combout ;
wire \ex_csr_addr[2]~q ;
wire \io_sw_r_ex_imm[2]~5_combout ;
wire \io_sw_r_ex_imm[2]~6_combout ;
wire \mem_imm~17_combout ;
wire \mem_imm[2]~q ;
wire \_T_3862[2]~4_combout ;
wire \pc_cntr[19]~7_combout ;
wire \pc_cntr[19]~8_combout ;
wire \npc[2]~0_combout ;
wire \pc_cntr~9_combout ;
wire \pc_cntr~10_combout ;
wire \pc_cntr~11_combout ;
wire \pc_cntr[19]~12_combout ;
wire \pc_cntr[2]~q ;
wire \id_pc~1_combout ;
wire \ex_pc~5_combout ;
wire \ex_pc[3]~q ;
wire \mem_pc~1_combout ;
wire \mem_pc[3]~q ;
wire \ex_inst~8_combout ;
wire \ex_inst[10]~q ;
wire \ex_inst~3_combout ;
wire \ex_inst[18]~q ;
wire \ex_csr_addr~3_combout ;
wire \ex_csr_addr[3]~q ;
wire \io_sw_r_ex_imm[3]~7_combout ;
wire \io_sw_r_ex_imm[3]~8_combout ;
wire \mem_imm~18_combout ;
wire \mem_imm[3]~q ;
wire \_T_3862[2]~5 ;
wire \_T_3862[3]~6_combout ;
wire \npc[2]~1 ;
wire \npc[3]~2_combout ;
wire \pc_cntr~13_combout ;
wire \pc_cntr~14_combout ;
wire \pc_cntr~15_combout ;
wire \pc_cntr[3]~q ;
wire \id_pc~2_combout ;
wire \ex_pc~0_combout ;
wire \ex_pc[4]~q ;
wire \mem_pc~2_combout ;
wire \mem_pc[4]~q ;
wire \ex_inst~9_combout ;
wire \ex_inst[11]~q ;
wire \ex_inst~4_combout ;
wire \ex_inst[19]~q ;
wire \ex_csr_addr~4_combout ;
wire \ex_csr_addr[4]~q ;
wire \io_sw_r_ex_imm[4]~3_combout ;
wire \io_sw_r_ex_imm[4]~4_combout ;
wire \mem_imm~19_combout ;
wire \mem_imm[4]~q ;
wire \_T_3862[3]~7 ;
wire \_T_3862[4]~8_combout ;
wire \ex_ctrl_alu_op2~6_combout ;
wire \ex_ctrl_alu_op2~7_combout ;
wire \ex_ctrl_alu_op2.01~q ;
wire \ex_ctrl_alu_op2~8_combout ;
wire \ex_ctrl_alu_op2.10~q ;
wire \csr_io_alu_op2[1]~0_combout ;
wire \ex_csr_cmd~4_combout ;
wire \ex_ctrl_alu_func~5_combout ;
wire \ex_ctrl_csr_cmd~11_combout ;
wire \Equal45~0_combout ;
wire \ex_ctrl_csr_cmd~12_combout ;
wire \Equal48~4_combout ;
wire \ex_ctrl_wb_sel~10_combout ;
wire \Equal50~0_combout ;
wire \ex_ctrl_csr_cmd~13_combout ;
wire \Equal51~0_combout ;
wire \ex_ctrl_csr_cmd~16_combout ;
wire \ex_ctrl_csr_cmd.000~q ;
wire \mem_ctrl_csr_cmd~14_combout ;
wire \mem_ctrl_csr_cmd.000~q ;
wire \mem_reg_waddr~1_combout ;
wire \mem_reg_waddr[1]~q ;
wire \mem_reg_waddr~0_combout ;
wire \mem_reg_waddr[0]~q ;
wire \_T_3681~0_combout ;
wire \mem_reg_waddr~3_combout ;
wire \mem_reg_waddr[3]~q ;
wire \mem_reg_waddr~2_combout ;
wire \mem_reg_waddr[2]~q ;
wire \_T_3681~1_combout ;
wire \_T_3681~2_combout ;
wire \mem_reg_waddr~4_combout ;
wire \mem_reg_waddr[4]~q ;
wire \Equal63~0_combout ;
wire \Equal62~0_combout ;
wire \Equal62~1_combout ;
wire \_T_3681~3_combout ;
wire \mem_csr_data~25_combout ;
wire \mem_csr_data[4]~q ;
wire \ex_ctrl_rf_wen~0_combout ;
wire \ex_ctrl_alu_op1~4_combout ;
wire \ex_ctrl_alu_op1~5_combout ;
wire \ex_ctrl_rf_wen~1_combout ;
wire \ex_ctrl_rf_wen~q ;
wire \mem_ctrl_rf_wen~0_combout ;
wire \mem_ctrl_rf_wen~q ;
wire \_T_3686~0_combout ;
wire \ex_rs_1[23]~0_combout ;
wire \ex_rs_1[23]~1_combout ;
wire \wb_ctrl_rf_wen~0_combout ;
wire \wb_ctrl_rf_wen~q ;
wire \wb_reg_waddr~4_combout ;
wire \wb_reg_waddr[4]~q ;
wire \wb_reg_waddr~0_combout ;
wire \wb_reg_waddr[0]~q ;
wire \wb_reg_waddr~1_combout ;
wire \wb_reg_waddr[1]~q ;
wire \wb_reg_waddr~2_combout ;
wire \wb_reg_waddr[2]~q ;
wire \wb_reg_waddr~3_combout ;
wire \wb_reg_waddr[3]~q ;
wire \_T_3543__T_3854_en~0_combout ;
wire \_T_3543__T_3854_en~1_combout ;
wire \wb_csr_data~18_combout ;
wire \wb_csr_data[4]~q ;
wire \wb_ctrl_wb_sel~14_combout ;
wire \wb_ctrl_wb_sel.10~q ;
wire \ex_ctrl_wb_sel~11_combout ;
wire \ex_ctrl_wb_sel~18_combout ;
wire \ex_ctrl_wb_sel~19_combout ;
wire \ex_ctrl_wb_sel.11~q ;
wire \mem_ctrl_wb_sel~13_combout ;
wire \mem_ctrl_wb_sel.11~q ;
wire \wb_ctrl_wb_sel~13_combout ;
wire \wb_ctrl_wb_sel.11~q ;
wire \_T_3543__T_3854_data[23]~2_combout ;
wire \npc[3]~3 ;
wire \npc[4]~4_combout ;
wire \id_npc~18_combout ;
wire \id_npc[4]~q ;
wire \ex_npc~18_combout ;
wire \ex_npc[4]~q ;
wire \mem_npc~16_combout ;
wire \mem_npc[4]~q ;
wire \wb_npc~16_combout ;
wire \wb_npc[4]~q ;
wire \ex_ctrl_wb_sel~13_combout ;
wire \ex_ctrl_wb_sel~14_combout ;
wire \ex_ctrl_wb_sel~15_combout ;
wire \ex_ctrl_wb_sel~12_combout ;
wire \ex_ctrl_wb_sel~16_combout ;
wire \ex_ctrl_wb_sel~17_combout ;
wire \ex_ctrl_wb_sel.00~q ;
wire \mem_ctrl_wb_sel~12_combout ;
wire \mem_ctrl_wb_sel.00~q ;
wire \wb_ctrl_wb_sel~12_combout ;
wire \wb_ctrl_wb_sel.00~q ;
wire \_T_3543__T_3854_data[23]~1_combout ;
wire \wb_alu_out~18_combout ;
wire \wb_alu_out[4]~q ;
wire \_T_3543__T_3854_data[4]~39_combout ;
wire \wb_dmem_read_data~60_combout ;
wire \ex_ctrl_mask_type~4_combout ;
wire \ex_ctrl_mask_type~5_combout ;
wire \ex_ctrl_mask_type~6_combout ;
wire \ex_ctrl_mask_type[0]~q ;
wire \mem_ctrl_mask_type~0_combout ;
wire \mem_ctrl_mask_type[0]~q ;
wire \ex_ctrl_mask_type~8_combout ;
wire \ex_ctrl_mask_type~9_combout ;
wire \ex_ctrl_mask_type~10_combout ;
wire \ex_ctrl_mask_type[1]~q ;
wire \mem_ctrl_mask_type~2_combout ;
wire \mem_ctrl_mask_type[1]~q ;
wire \wb_dmem_read_data[7]~17_combout ;
wire \wb_dmem_read_data[4]~4_combout ;
wire \wb_dmem_read_data[7]~18_combout ;
wire \wb_dmem_read_data[7]~19_combout ;
wire \wb_dmem_read_data[7]~20_combout ;
wire \wb_dmem_read_data[7]~21_combout ;
wire \wb_dmem_read_data[4]~q ;
wire \_T_3543__T_3854_data[4]~40_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a28~portbdataout ;
wire \ex_rs_1~20_combout ;
wire \ex_rs_1[4]~q ;
wire \wb_ctrl_csr_cmd~14_combout ;
wire \wb_ctrl_csr_cmd.000~q ;
wire \Equal53~1_combout ;
wire \_T_3091~combout ;
wire \_GEN_15~combout ;
wire \ex_ctrl_mem_en~q ;
wire \ex_reg_rs1_bypass[2]~8_combout ;
wire \Equal64~0_combout ;
wire \_T_3689~0_combout ;
wire \_T_3689~1_combout ;
wire \_T_3689~2_combout ;
wire \ex_reg_rs2_bypass[7]~4_combout ;
wire \_GEN_39~combout ;
wire \mem_ctrl_mem_en~q ;
wire \wb_ctrl_mem_en~0_combout ;
wire \wb_ctrl_mem_en~q ;
wire \ex_reg_rs1_bypass[2]~6_combout ;
wire \ex_reg_rs1_bypass[2]~12_combout ;
wire \ex_reg_rs2_bypass[7]~5_combout ;
wire \ex_reg_rs2_bypass[4]~75_combout ;
wire \ex_reg_rs2_bypass[4]~76_combout ;
wire \alu_io_op2[4]~60_combout ;
wire \alu_io_op2[4]~61_combout ;
wire \alu_io_op2[4]~62_combout ;
wire \ex_ctrl_alu_func~16_combout ;
wire \Equal35~0_combout ;
wire \Equal36~0_combout ;
wire \ex_ctrl_alu_func~17_combout ;
wire \ex_ctrl_alu_func~18_combout ;
wire \ex_ctrl_alu_func~19_combout ;
wire \ex_ctrl_alu_func~20_combout ;
wire \ex_ctrl_alu_func~21_combout ;
wire \ex_ctrl_alu_func~22_combout ;
wire \ex_ctrl_alu_func~23_combout ;
wire \ex_ctrl_alu_func[3]~q ;
wire \ex_ctrl_alu_func~24_combout ;
wire \ex_ctrl_alu_func~25_combout ;
wire \ex_ctrl_alu_func~26_combout ;
wire \ex_ctrl_alu_func~27_combout ;
wire \ex_ctrl_alu_func~35_combout ;
wire \ex_ctrl_alu_func~36_combout ;
wire \ex_ctrl_alu_func~28_combout ;
wire \ex_ctrl_alu_func[1]~q ;
wire \ex_ctrl_alu_func~29_combout ;
wire \ex_ctrl_alu_func~30_combout ;
wire \ex_ctrl_alu_func~31_combout ;
wire \ex_ctrl_alu_func~32_combout ;
wire \ex_ctrl_alu_func[2]~q ;
wire \mem_alu_out[26]~0_combout ;
wire \ex_ctrl_alu_op1~6_combout ;
wire \ex_ctrl_alu_op1[0]~q ;
wire \ex_ctrl_alu_op1[1]~q ;
wire \Equal59~0_combout ;
wire \Equal59~1_combout ;
wire \Equal60~2_combout ;
wire \Equal60~3_combout ;
wire \Equal60~5_combout ;
wire \Equal60~4_combout ;
wire \csr_io_in[0]~0_combout ;
wire \ex_reg_rs1_bypass[0]~4_combout ;
wire \ex_reg_rs1_bypass[0]~20_combout ;
wire \_T_3634~2_combout ;
wire \ex_reg_rs1_bypass[4]~82_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a28~portbdataout ;
wire \ex_rs_0~20_combout ;
wire \ex_rs_0[4]~q ;
wire \Equal61~0_combout ;
wire \Equal61~1_combout ;
wire \Equal61~2_combout ;
wire \ex_reg_rs1_bypass[2]~138_combout ;
wire \ex_reg_rs1_bypass[2]~7_combout ;
wire \ex_reg_rs1_bypass[4]~83_combout ;
wire \ex_reg_rs1_bypass[4]~84_combout ;
wire \ex_reg_rs1_bypass[4]~85_combout ;
wire \alu_io_op1[4]~106_combout ;
wire \mem_alu_out[26]~1_combout ;
wire \mem_alu_out[26]~2_combout ;
wire \mem_alu_out~143_combout ;
wire \mem_alu_out~144_combout ;
wire \mem_alu_out~85_combout ;
wire \mem_alu_out~86_combout ;
wire \mem_alu_out[26]~5_combout ;
wire \mem_alu_out[26]~6_combout ;
wire \mem_alu_out~87_combout ;
wire \mem_alu_out[4]~q ;
wire \pc_cntr~16_combout ;
wire \pc_cntr~17_combout ;
wire \pc_cntr~18_combout ;
wire \pc_cntr[4]~q ;
wire \id_pc~3_combout ;
wire \ex_pc~1_combout ;
wire \ex_pc[5]~q ;
wire \mem_csr_data~28_combout ;
wire \mem_csr_data[5]~q ;
wire \ex_reg_rs1_bypass[5]~90_combout ;
wire \wb_csr_data~21_combout ;
wire \wb_csr_data[5]~q ;
wire \npc[4]~5 ;
wire \npc[5]~6_combout ;
wire \id_npc~21_combout ;
wire \id_npc[5]~q ;
wire \ex_npc~21_combout ;
wire \ex_npc[5]~q ;
wire \mem_npc~19_combout ;
wire \mem_npc[5]~q ;
wire \wb_npc~19_combout ;
wire \wb_npc[5]~q ;
wire \wb_alu_out~21_combout ;
wire \wb_alu_out[5]~q ;
wire \_T_3543__T_3854_data[5]~45_combout ;
wire \wb_dmem_read_data~64_combout ;
wire \wb_dmem_read_data[5]~3_combout ;
wire \wb_dmem_read_data[5]~q ;
wire \_T_3543__T_3854_data[5]~46_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a27~portbdataout ;
wire \ex_rs_0~22_combout ;
wire \ex_rs_0[5]~q ;
wire \ex_reg_rs1_bypass[5]~91_combout ;
wire \ex_reg_rs1_bypass[5]~92_combout ;
wire \ex_reg_rs1_bypass[5]~93_combout ;
wire \alu_io_op1[5]~108_combout ;
wire \alu_io_op2[5]~43_combout ;
wire \ex_csr_addr~9_combout ;
wire \ex_csr_addr[5]~q ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a27~portbdataout ;
wire \ex_rs_1~23_combout ;
wire \ex_rs_1[5]~q ;
wire \ex_reg_rs2_bypass[5]~83_combout ;
wire \ex_reg_rs2_bypass[5]~84_combout ;
wire \ex_reg_rs2_bypass[5]~85_combout ;
wire \alu_io_op2[5]~67_combout ;
wire \alu_io_op2[5]~68_combout ;
wire \mem_alu_out~141_combout ;
wire \mem_alu_out~142_combout ;
wire \mem_alu_out~88_combout ;
wire \mem_alu_out~89_combout ;
wire \mem_alu_out~90_combout ;
wire \mem_alu_out[5]~q ;
wire \mem_pc~3_combout ;
wire \mem_pc[5]~q ;
wire \mem_imm~20_combout ;
wire \mem_imm[5]~q ;
wire \_T_3862[4]~9 ;
wire \_T_3862[5]~10_combout ;
wire \pc_cntr~19_combout ;
wire \pc_cntr~20_combout ;
wire \pc_cntr~21_combout ;
wire \pc_cntr[5]~q ;
wire \id_pc~4_combout ;
wire \ex_pc~2_combout ;
wire \ex_pc[6]~q ;
wire \mem_pc~4_combout ;
wire \mem_pc[6]~q ;
wire \ex_csr_addr~10_combout ;
wire \ex_csr_addr[6]~q ;
wire \mem_imm~21_combout ;
wire \mem_imm[6]~q ;
wire \_T_3862[5]~11 ;
wire \_T_3862[6]~12_combout ;
wire \mem_csr_data~29_combout ;
wire \mem_csr_data[6]~q ;
wire \wb_csr_data~22_combout ;
wire \wb_csr_data[6]~q ;
wire \npc[5]~7 ;
wire \npc[6]~8_combout ;
wire \id_npc~22_combout ;
wire \id_npc[6]~q ;
wire \ex_npc~22_combout ;
wire \ex_npc[6]~q ;
wire \mem_npc~20_combout ;
wire \mem_npc[6]~q ;
wire \wb_npc~20_combout ;
wire \wb_npc[6]~q ;
wire \wb_alu_out~22_combout ;
wire \wb_alu_out[6]~q ;
wire \_T_3543__T_3854_data[6]~47_combout ;
wire \wb_dmem_read_data~68_combout ;
wire \wb_dmem_read_data[6]~2_combout ;
wire \wb_dmem_read_data[6]~q ;
wire \_T_3543__T_3854_data[6]~48_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a26~portbdataout ;
wire \ex_rs_1~24_combout ;
wire \ex_rs_1[6]~q ;
wire \ex_reg_rs2_bypass[6]~86_combout ;
wire \ex_reg_rs2_bypass[6]~87_combout ;
wire \ex_reg_rs2_bypass[6]~88_combout ;
wire \alu_io_op2[6]~69_combout ;
wire \alu_io_op2[6]~70_combout ;
wire \ex_reg_rs1_bypass[6]~98_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a26~portbdataout ;
wire \ex_rs_0~24_combout ;
wire \ex_rs_0[6]~q ;
wire \ex_reg_rs1_bypass[6]~99_combout ;
wire \ex_reg_rs1_bypass[6]~100_combout ;
wire \ex_reg_rs1_bypass[6]~101_combout ;
wire \alu_io_op1[6]~110_combout ;
wire \mem_alu_out~139_combout ;
wire \mem_alu_out~140_combout ;
wire \mem_alu_out~91_combout ;
wire \mem_alu_out~92_combout ;
wire \mem_alu_out~93_combout ;
wire \mem_alu_out[6]~q ;
wire \pc_cntr~22_combout ;
wire \pc_cntr~23_combout ;
wire \pc_cntr~24_combout ;
wire \pc_cntr[6]~q ;
wire \id_pc~5_combout ;
wire \ex_pc~3_combout ;
wire \ex_pc[7]~q ;
wire \mem_csr_data~30_combout ;
wire \mem_csr_data[7]~q ;
wire \ex_reg_rs1_bypass[7]~102_combout ;
wire \wb_csr_data~23_combout ;
wire \wb_csr_data[7]~q ;
wire \npc[6]~9 ;
wire \npc[7]~10_combout ;
wire \id_npc~23_combout ;
wire \id_npc[7]~q ;
wire \ex_npc~23_combout ;
wire \ex_npc[7]~q ;
wire \mem_npc~21_combout ;
wire \mem_npc[7]~q ;
wire \wb_npc~21_combout ;
wire \wb_npc[7]~q ;
wire \wb_alu_out~23_combout ;
wire \wb_alu_out[7]~q ;
wire \_T_3543__T_3854_data[7]~49_combout ;
wire \wb_dmem_read_data~28_combout ;
wire \wb_dmem_read_data[7]~1_combout ;
wire \wb_dmem_read_data[7]~q ;
wire \_T_3543__T_3854_data[7]~50_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a25~portbdataout ;
wire \ex_rs_0~25_combout ;
wire \ex_rs_0[7]~q ;
wire \ex_reg_rs1_bypass[7]~103_combout ;
wire \ex_reg_rs1_bypass[7]~104_combout ;
wire \ex_reg_rs1_bypass[7]~105_combout ;
wire \alu_io_op1[7]~111_combout ;
wire \ex_csr_addr~11_combout ;
wire \ex_csr_addr[7]~q ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a25~portbdataout ;
wire \ex_rs_1~25_combout ;
wire \ex_rs_1[7]~q ;
wire \ex_reg_rs2_bypass[7]~89_combout ;
wire \ex_reg_rs2_bypass[7]~90_combout ;
wire \ex_reg_rs2_bypass[7]~91_combout ;
wire \alu_io_op2[7]~71_combout ;
wire \alu_io_op2[7]~72_combout ;
wire \mem_alu_out~94_combout ;
wire \mem_alu_out~95_combout ;
wire \mem_alu_out~96_combout ;
wire \mem_alu_out~97_combout ;
wire \mem_alu_out~98_combout ;
wire \mem_alu_out[7]~q ;
wire \mem_pc~5_combout ;
wire \mem_pc[7]~q ;
wire \mem_imm~22_combout ;
wire \mem_imm[7]~q ;
wire \_T_3862[6]~13 ;
wire \_T_3862[7]~14_combout ;
wire \pc_cntr~25_combout ;
wire \pc_cntr~26_combout ;
wire \pc_cntr~27_combout ;
wire \pc_cntr[7]~q ;
wire \id_pc~6_combout ;
wire \ex_pc~6_combout ;
wire \ex_pc[8]~q ;
wire \mem_pc~6_combout ;
wire \mem_pc[8]~q ;
wire \ex_csr_addr~5_combout ;
wire \ex_csr_addr[8]~q ;
wire \mem_imm~23_combout ;
wire \mem_imm[8]~q ;
wire \_T_3862[7]~15 ;
wire \_T_3862[8]~16_combout ;
wire \mem_csr_data~13_combout ;
wire \mem_csr_data[8]~q ;
wire \wb_csr_data~6_combout ;
wire \wb_csr_data[8]~q ;
wire \npc[7]~11 ;
wire \npc[8]~12_combout ;
wire \id_npc~6_combout ;
wire \id_npc[8]~q ;
wire \ex_npc~6_combout ;
wire \ex_npc[8]~q ;
wire \mem_npc~4_combout ;
wire \mem_npc[8]~q ;
wire \wb_npc~4_combout ;
wire \wb_npc[8]~q ;
wire \wb_alu_out~6_combout ;
wire \wb_alu_out[8]~q ;
wire \_T_3543__T_3854_data[8]~15_combout ;
wire \wb_dmem_read_data[22]~89_combout ;
wire \wb_dmem_read_data[22]~90_combout ;
wire \wb_dmem_read_data~22_combout ;
wire \wb_dmem_read_data~43_combout ;
wire \wb_dmem_read_data~44_combout ;
wire \wb_dmem_read_data[14]~45_combout ;
wire \wb_dmem_read_data[14]~46_combout ;
wire \wb_dmem_read_data[14]~47_combout ;
wire \wb_dmem_read_data~48_combout ;
wire \wb_dmem_read_data[8]~q ;
wire \_T_3543__T_3854_data[8]~16_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a24~portbdataout ;
wire \ex_rs_1~9_combout ;
wire \ex_rs_1[8]~q ;
wire \ex_reg_rs2_bypass[8]~34_combout ;
wire \ex_reg_rs2_bypass[8]~35_combout ;
wire \ex_reg_rs2_bypass[8]~36_combout ;
wire \alu_io_op2[8]~46_combout ;
wire \alu_io_op2[8]~47_combout ;
wire \ex_reg_rs1_bypass[8]~34_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a24~portbdataout ;
wire \ex_rs_0~8_combout ;
wire \ex_rs_0[8]~q ;
wire \ex_reg_rs1_bypass[8]~35_combout ;
wire \ex_reg_rs1_bypass[8]~36_combout ;
wire \ex_reg_rs1_bypass[8]~37_combout ;
wire \alu_io_op1[8]~94_combout ;
wire \mem_alu_out~155_combout ;
wire \mem_alu_out~156_combout ;
wire \mem_alu_out~37_combout ;
wire \mem_alu_out~38_combout ;
wire \mem_alu_out~39_combout ;
wire \mem_alu_out[8]~q ;
wire \pc_cntr~28_combout ;
wire \pc_cntr~29_combout ;
wire \pc_cntr~30_combout ;
wire \pc_cntr[8]~q ;
wire \id_pc~7_combout ;
wire \ex_pc~7_combout ;
wire \ex_pc[9]~q ;
wire \mem_csr_data~14_combout ;
wire \mem_csr_data[9]~q ;
wire \ex_reg_rs1_bypass[9]~38_combout ;
wire \wb_csr_data~7_combout ;
wire \wb_csr_data[9]~q ;
wire \npc[8]~13 ;
wire \npc[9]~14_combout ;
wire \id_npc~7_combout ;
wire \id_npc[9]~q ;
wire \ex_npc~7_combout ;
wire \ex_npc[9]~q ;
wire \mem_npc~5_combout ;
wire \mem_npc[9]~q ;
wire \wb_npc~5_combout ;
wire \wb_npc[9]~q ;
wire \wb_alu_out~7_combout ;
wire \wb_alu_out[9]~q ;
wire \_T_3543__T_3854_data[9]~17_combout ;
wire \wb_dmem_read_data~16_combout ;
wire \wb_dmem_read_data~49_combout ;
wire \wb_dmem_read_data~50_combout ;
wire \wb_dmem_read_data~51_combout ;
wire \wb_dmem_read_data[9]~q ;
wire \_T_3543__T_3854_data[9]~18_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a23~portbdataout ;
wire \ex_rs_0~9_combout ;
wire \ex_rs_0[9]~q ;
wire \ex_reg_rs1_bypass[9]~39_combout ;
wire \ex_reg_rs1_bypass[9]~40_combout ;
wire \ex_reg_rs1_bypass[9]~41_combout ;
wire \alu_io_op1[9]~95_combout ;
wire \ex_csr_addr~6_combout ;
wire \ex_csr_addr[9]~q ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a23~portbdataout ;
wire \ex_rs_1~8_combout ;
wire \ex_rs_1[9]~q ;
wire \ex_reg_rs2_bypass[9]~31_combout ;
wire \ex_reg_rs2_bypass[9]~32_combout ;
wire \ex_reg_rs2_bypass[9]~33_combout ;
wire \alu_io_op2[9]~44_combout ;
wire \alu_io_op2[9]~45_combout ;
wire \mem_alu_out~153_combout ;
wire \mem_alu_out~154_combout ;
wire \mem_alu_out~40_combout ;
wire \mem_alu_out~41_combout ;
wire \mem_alu_out~42_combout ;
wire \mem_alu_out[9]~q ;
wire \mem_pc~7_combout ;
wire \mem_pc[9]~q ;
wire \mem_imm~24_combout ;
wire \mem_imm[9]~q ;
wire \_T_3862[8]~17 ;
wire \_T_3862[9]~18_combout ;
wire \pc_cntr~31_combout ;
wire \pc_cntr~32_combout ;
wire \pc_cntr~33_combout ;
wire \pc_cntr[9]~q ;
wire \id_pc~8_combout ;
wire \ex_pc~8_combout ;
wire \ex_pc[10]~q ;
wire \mem_pc~8_combout ;
wire \mem_pc[10]~q ;
wire \ex_csr_addr~8_combout ;
wire \ex_csr_addr[10]~q ;
wire \mem_imm~25_combout ;
wire \mem_imm[10]~q ;
wire \_T_3862[9]~19 ;
wire \_T_3862[10]~20_combout ;
wire \mem_csr_data~15_combout ;
wire \mem_csr_data[10]~q ;
wire \wb_csr_data~8_combout ;
wire \wb_csr_data[10]~q ;
wire \npc[9]~15 ;
wire \npc[10]~16_combout ;
wire \id_npc~8_combout ;
wire \id_npc[10]~q ;
wire \ex_npc~8_combout ;
wire \ex_npc[10]~q ;
wire \mem_npc~6_combout ;
wire \mem_npc[10]~q ;
wire \wb_npc~6_combout ;
wire \wb_npc[10]~q ;
wire \wb_alu_out~8_combout ;
wire \wb_alu_out[10]~q ;
wire \_T_3543__T_3854_data[10]~19_combout ;
wire \wb_dmem_read_data~52_combout ;
wire \wb_dmem_read_data~53_combout ;
wire \wb_dmem_read_data~54_combout ;
wire \wb_dmem_read_data~55_combout ;
wire \wb_dmem_read_data[10]~q ;
wire \_T_3543__T_3854_data[10]~20_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a22~portbdataout ;
wire \ex_rs_1~10_combout ;
wire \ex_rs_1[10]~q ;
wire \ex_reg_rs2_bypass[10]~37_combout ;
wire \ex_reg_rs2_bypass[10]~38_combout ;
wire \ex_reg_rs2_bypass[10]~39_combout ;
wire \alu_io_op2[10]~48_combout ;
wire \alu_io_op2[10]~49_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a22~portbdataout ;
wire \ex_rs_0~10_combout ;
wire \ex_rs_0[10]~q ;
wire \ex_reg_rs1_bypass[10]~42_combout ;
wire \ex_reg_rs1_bypass[10]~43_combout ;
wire \ex_reg_rs1_bypass[10]~44_combout ;
wire \ex_reg_rs1_bypass[10]~139_combout ;
wire \ex_reg_rs1_bypass[10]~45_combout ;
wire \alu_io_op1[10]~96_combout ;
wire \mem_alu_out~151_combout ;
wire \mem_alu_out~152_combout ;
wire \mem_alu_out~43_combout ;
wire \mem_alu_out~44_combout ;
wire \mem_alu_out~45_combout ;
wire \mem_alu_out[10]~q ;
wire \pc_cntr~34_combout ;
wire \pc_cntr~35_combout ;
wire \pc_cntr~36_combout ;
wire \pc_cntr[10]~q ;
wire \id_pc~9_combout ;
wire \ex_pc~9_combout ;
wire \ex_pc[11]~q ;
wire \mem_csr_data~16_combout ;
wire \mem_csr_data[11]~q ;
wire \ex_reg_rs1_bypass[11]~46_combout ;
wire \wb_csr_data~9_combout ;
wire \wb_csr_data[11]~q ;
wire \npc[10]~17 ;
wire \npc[11]~18_combout ;
wire \id_npc~9_combout ;
wire \id_npc[11]~q ;
wire \ex_npc~9_combout ;
wire \ex_npc[11]~q ;
wire \mem_npc~7_combout ;
wire \mem_npc[11]~q ;
wire \wb_npc~7_combout ;
wire \wb_npc[11]~q ;
wire \wb_alu_out~9_combout ;
wire \wb_alu_out[11]~q ;
wire \_T_3543__T_3854_data[11]~21_combout ;
wire \wb_dmem_read_data~56_combout ;
wire \wb_dmem_read_data~57_combout ;
wire \wb_dmem_read_data~58_combout ;
wire \wb_dmem_read_data~59_combout ;
wire \wb_dmem_read_data[11]~q ;
wire \_T_3543__T_3854_data[11]~22_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a21~portbdataout ;
wire \ex_rs_0~11_combout ;
wire \ex_rs_0[11]~q ;
wire \ex_reg_rs1_bypass[11]~47_combout ;
wire \ex_reg_rs1_bypass[11]~48_combout ;
wire \ex_reg_rs1_bypass[11]~49_combout ;
wire \alu_io_op1[11]~97_combout ;
wire \ex_csr_addr~7_combout ;
wire \ex_csr_addr[11]~q ;
wire \_T_3593~0_combout ;
wire \ex_ctrl_imm_type~21_combout ;
wire \ex_ctrl_imm_type.100~q ;
wire \_T_3593~1_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a21~portbdataout ;
wire \ex_rs_1~11_combout ;
wire \ex_rs_1[11]~q ;
wire \ex_reg_rs2_bypass[11]~40_combout ;
wire \ex_reg_rs2_bypass[11]~41_combout ;
wire \ex_reg_rs2_bypass[11]~42_combout ;
wire \alu_io_op2[11]~50_combout ;
wire \alu_io_op2[11]~51_combout ;
wire \mem_alu_out~46_combout ;
wire \mem_alu_out~47_combout ;
wire \mem_alu_out~48_combout ;
wire \mem_alu_out~49_combout ;
wire \mem_alu_out~50_combout ;
wire \mem_alu_out[11]~q ;
wire \mem_pc~9_combout ;
wire \mem_pc[11]~q ;
wire \mem_imm~26_combout ;
wire \mem_imm[11]~q ;
wire \_T_3862[10]~21 ;
wire \_T_3862[11]~22_combout ;
wire \pc_cntr~37_combout ;
wire \pc_cntr~38_combout ;
wire \pc_cntr~39_combout ;
wire \pc_cntr[11]~q ;
wire \id_pc~10_combout ;
wire \ex_pc~10_combout ;
wire \ex_pc[12]~q ;
wire \mem_pc~10_combout ;
wire \mem_pc[12]~q ;
wire \ex_inst~11_combout ;
wire \ex_inst[12]~q ;
wire \mem_imm~7_combout ;
wire \_T_3579~combout ;
wire \mem_imm~27_combout ;
wire \mem_imm[12]~q ;
wire \_T_3862[11]~23 ;
wire \_T_3862[12]~24_combout ;
wire \alu_io_op2[12]~53_combout ;
wire \mem_csr_data~17_combout ;
wire \mem_csr_data[12]~q ;
wire \wb_csr_data~10_combout ;
wire \wb_csr_data[12]~q ;
wire \npc[11]~19 ;
wire \npc[12]~20_combout ;
wire \id_npc~10_combout ;
wire \id_npc[12]~q ;
wire \ex_npc~10_combout ;
wire \ex_npc[12]~q ;
wire \mem_npc~8_combout ;
wire \mem_npc[12]~q ;
wire \wb_npc~8_combout ;
wire \wb_npc[12]~q ;
wire \wb_alu_out~10_combout ;
wire \wb_alu_out[12]~q ;
wire \_T_3543__T_3854_data[12]~23_combout ;
wire \wb_dmem_read_data~61_combout ;
wire \wb_dmem_read_data~62_combout ;
wire \wb_dmem_read_data~63_combout ;
wire \wb_dmem_read_data[12]~q ;
wire \_T_3543__T_3854_data[12]~24_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a20~portbdataout ;
wire \ex_rs_1~13_combout ;
wire \ex_rs_1[12]~q ;
wire \ex_reg_rs2_bypass[12]~47_combout ;
wire \ex_reg_rs2_bypass[12]~48_combout ;
wire \ex_reg_rs2_bypass[12]~49_combout ;
wire \ex_reg_rs2_bypass[12]~50_combout ;
wire \alu_io_op2[12]~78_combout ;
wire \ex_reg_rs1_bypass[12]~50_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a20~portbdataout ;
wire \ex_rs_0~12_combout ;
wire \ex_rs_0[12]~q ;
wire \ex_reg_rs1_bypass[12]~51_combout ;
wire \ex_reg_rs1_bypass[12]~52_combout ;
wire \ex_reg_rs1_bypass[12]~53_combout ;
wire \alu_io_op1[12]~98_combout ;
wire \mem_alu_out~149_combout ;
wire \mem_alu_out~150_combout ;
wire \mem_alu_out~51_combout ;
wire \mem_alu_out~52_combout ;
wire \mem_alu_out~53_combout ;
wire \mem_alu_out[12]~q ;
wire \pc_cntr~40_combout ;
wire \pc_cntr~41_combout ;
wire \pc_cntr~42_combout ;
wire \pc_cntr[12]~q ;
wire \id_pc~11_combout ;
wire \ex_pc~11_combout ;
wire \ex_pc[13]~q ;
wire \mem_csr_data~18_combout ;
wire \mem_csr_data[13]~q ;
wire \ex_reg_rs1_bypass[13]~54_combout ;
wire \wb_csr_data~11_combout ;
wire \wb_csr_data[13]~q ;
wire \npc[12]~21 ;
wire \npc[13]~22_combout ;
wire \id_npc~11_combout ;
wire \id_npc[13]~q ;
wire \ex_npc~11_combout ;
wire \ex_npc[13]~q ;
wire \mem_npc~9_combout ;
wire \mem_npc[13]~q ;
wire \wb_npc~9_combout ;
wire \wb_npc[13]~q ;
wire \wb_alu_out~11_combout ;
wire \wb_alu_out[13]~q ;
wire \_T_3543__T_3854_data[13]~25_combout ;
wire \wb_dmem_read_data~65_combout ;
wire \wb_dmem_read_data~66_combout ;
wire \wb_dmem_read_data~67_combout ;
wire \wb_dmem_read_data[13]~q ;
wire \_T_3543__T_3854_data[13]~26_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a19~portbdataout ;
wire \ex_rs_0~13_combout ;
wire \ex_rs_0[13]~q ;
wire \ex_reg_rs1_bypass[13]~55_combout ;
wire \ex_reg_rs1_bypass[13]~56_combout ;
wire \ex_reg_rs1_bypass[13]~57_combout ;
wire \alu_io_op1[13]~99_combout ;
wire \ex_inst~10_combout ;
wire \ex_inst[13]~q ;
wire \alu_io_op2[13]~52_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a19~portbdataout ;
wire \ex_rs_1~12_combout ;
wire \ex_rs_1[13]~q ;
wire \ex_reg_rs2_bypass[13]~43_combout ;
wire \ex_reg_rs2_bypass[13]~44_combout ;
wire \ex_reg_rs2_bypass[13]~45_combout ;
wire \ex_reg_rs2_bypass[13]~46_combout ;
wire \alu_io_op2[13]~77_combout ;
wire \mem_alu_out~54_combout ;
wire \mem_alu_out~55_combout ;
wire \mem_alu_out~56_combout ;
wire \mem_alu_out~57_combout ;
wire \mem_alu_out~58_combout ;
wire \mem_alu_out[13]~q ;
wire \mem_pc~11_combout ;
wire \mem_pc[13]~q ;
wire \mem_imm~28_combout ;
wire \mem_imm[13]~q ;
wire \_T_3862[12]~25 ;
wire \_T_3862[13]~26_combout ;
wire \pc_cntr~43_combout ;
wire \pc_cntr~44_combout ;
wire \pc_cntr~45_combout ;
wire \pc_cntr[13]~q ;
wire \id_pc~12_combout ;
wire \ex_pc~12_combout ;
wire \ex_pc[14]~q ;
wire \mem_pc~12_combout ;
wire \mem_pc[14]~q ;
wire \ex_inst~12_combout ;
wire \ex_inst[14]~q ;
wire \mem_imm~29_combout ;
wire \mem_imm[14]~q ;
wire \_T_3862[13]~27 ;
wire \_T_3862[14]~28_combout ;
wire \alu_io_op2[14]~54_combout ;
wire \mem_csr_data~19_combout ;
wire \mem_csr_data[14]~q ;
wire \wb_csr_data~12_combout ;
wire \wb_csr_data[14]~q ;
wire \npc[13]~23 ;
wire \npc[14]~24_combout ;
wire \id_npc~12_combout ;
wire \id_npc[14]~q ;
wire \ex_npc~12_combout ;
wire \ex_npc[14]~q ;
wire \mem_npc~10_combout ;
wire \mem_npc[14]~q ;
wire \wb_npc~10_combout ;
wire \wb_npc[14]~q ;
wire \wb_alu_out~12_combout ;
wire \wb_alu_out[14]~q ;
wire \_T_3543__T_3854_data[14]~27_combout ;
wire \wb_dmem_read_data~69_combout ;
wire \wb_dmem_read_data~70_combout ;
wire \wb_dmem_read_data~71_combout ;
wire \wb_dmem_read_data[14]~q ;
wire \_T_3543__T_3854_data[14]~28_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a18~portbdataout ;
wire \ex_rs_1~14_combout ;
wire \ex_rs_1[14]~q ;
wire \ex_reg_rs2_bypass[14]~51_combout ;
wire \ex_reg_rs2_bypass[14]~52_combout ;
wire \ex_reg_rs2_bypass[14]~53_combout ;
wire \ex_reg_rs2_bypass[14]~54_combout ;
wire \alu_io_op2[14]~79_combout ;
wire \ex_reg_rs1_bypass[14]~58_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a18~portbdataout ;
wire \ex_rs_0~14_combout ;
wire \ex_rs_0[14]~q ;
wire \ex_reg_rs1_bypass[14]~59_combout ;
wire \ex_reg_rs1_bypass[14]~60_combout ;
wire \ex_reg_rs1_bypass[14]~61_combout ;
wire \alu_io_op1[14]~100_combout ;
wire \mem_alu_out~147_combout ;
wire \mem_alu_out~148_combout ;
wire \mem_alu_out~59_combout ;
wire \mem_alu_out~60_combout ;
wire \mem_alu_out~61_combout ;
wire \mem_alu_out[14]~q ;
wire \pc_cntr~46_combout ;
wire \pc_cntr~47_combout ;
wire \pc_cntr~48_combout ;
wire \pc_cntr[14]~q ;
wire \id_pc~13_combout ;
wire \ex_pc~13_combout ;
wire \ex_pc[15]~q ;
wire \mem_csr_data~20_combout ;
wire \mem_csr_data[15]~q ;
wire \ex_reg_rs1_bypass[15]~62_combout ;
wire \wb_csr_data~13_combout ;
wire \wb_csr_data[15]~q ;
wire \npc[14]~25 ;
wire \npc[15]~26_combout ;
wire \id_npc~13_combout ;
wire \id_npc[15]~q ;
wire \ex_npc~13_combout ;
wire \ex_npc[15]~q ;
wire \mem_npc~11_combout ;
wire \mem_npc[15]~q ;
wire \wb_npc~11_combout ;
wire \wb_npc[15]~q ;
wire \wb_alu_out~13_combout ;
wire \wb_alu_out[15]~q ;
wire \_T_3543__T_3854_data[15]~29_combout ;
wire \wb_dmem_read_data~72_combout ;
wire \wb_dmem_read_data~91_combout ;
wire \Equal69~0_combout ;
wire \wb_dmem_read_data~39_combout ;
wire \wb_dmem_read_data~73_combout ;
wire \wb_dmem_read_data~74_combout ;
wire \wb_dmem_read_data[15]~q ;
wire \_T_3543__T_3854_data[15]~30_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a17~portbdataout ;
wire \ex_rs_0~15_combout ;
wire \ex_rs_0[15]~q ;
wire \ex_reg_rs1_bypass[15]~63_combout ;
wire \ex_reg_rs1_bypass[15]~64_combout ;
wire \ex_reg_rs1_bypass[15]~65_combout ;
wire \alu_io_op1[15]~101_combout ;
wire \alu_io_op2[15]~55_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a17~portbdataout ;
wire \ex_rs_1~15_combout ;
wire \ex_rs_1[15]~q ;
wire \ex_reg_rs2_bypass[15]~55_combout ;
wire \ex_reg_rs2_bypass[15]~56_combout ;
wire \ex_reg_rs2_bypass[15]~57_combout ;
wire \ex_reg_rs2_bypass[15]~58_combout ;
wire \alu_io_op2[15]~92_combout ;
wire \mem_alu_out~62_combout ;
wire \mem_alu_out~63_combout ;
wire \mem_alu_out~64_combout ;
wire \mem_alu_out~65_combout ;
wire \mem_alu_out~66_combout ;
wire \mem_alu_out[15]~q ;
wire \mem_pc~13_combout ;
wire \mem_pc[15]~q ;
wire \mem_imm~30_combout ;
wire \mem_imm[15]~q ;
wire \_T_3862[14]~29 ;
wire \_T_3862[15]~30_combout ;
wire \pc_cntr~49_combout ;
wire \pc_cntr~50_combout ;
wire \pc_cntr~51_combout ;
wire \pc_cntr[15]~q ;
wire \id_pc~14_combout ;
wire \ex_pc~14_combout ;
wire \ex_pc[16]~q ;
wire \mem_pc~14_combout ;
wire \mem_pc[16]~q ;
wire \mem_imm~31_combout ;
wire \mem_imm[16]~q ;
wire \_T_3862[15]~31 ;
wire \_T_3862[16]~32_combout ;
wire \alu_io_op2[16]~57_combout ;
wire \mem_csr_data~21_combout ;
wire \mem_csr_data[16]~q ;
wire \wb_csr_data~14_combout ;
wire \wb_csr_data[16]~q ;
wire \npc[15]~27 ;
wire \npc[16]~28_combout ;
wire \id_npc~14_combout ;
wire \id_npc[16]~q ;
wire \ex_npc~14_combout ;
wire \ex_npc[16]~q ;
wire \mem_npc~12_combout ;
wire \mem_npc[16]~q ;
wire \wb_npc~12_combout ;
wire \wb_npc[16]~q ;
wire \wb_alu_out~14_combout ;
wire \wb_alu_out[16]~q ;
wire \_T_3543__T_3854_data[16]~31_combout ;
wire \wb_dmem_read_data~23_combout ;
wire \ex_ctrl_wb_sel~20_combout ;
wire \ex_ctrl_mask_type~7_combout ;
wire \ex_ctrl_mask_type[2]~q ;
wire \mem_ctrl_mask_type~1_combout ;
wire \mem_ctrl_mask_type[2]~q ;
wire \wb_dmem_read_data[22]~24_combout ;
wire \wb_dmem_read_data[22]~25_combout ;
wire \wb_dmem_read_data~26_combout ;
wire \wb_dmem_read_data~34_combout ;
wire \wb_dmem_read_data~35_combout ;
wire \Equal68~1_combout ;
wire \wb_dmem_read_data~36_combout ;
wire \wb_dmem_read_data[22]~31_combout ;
wire \wb_dmem_read_data[22]~32_combout ;
wire \wb_dmem_read_data~75_combout ;
wire \wb_dmem_read_data[16]~q ;
wire \_T_3543__T_3854_data[16]~32_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a16~portbdataout ;
wire \ex_rs_1~17_combout ;
wire \ex_rs_1[16]~q ;
wire \ex_reg_rs2_bypass[16]~63_combout ;
wire \ex_reg_rs2_bypass[16]~64_combout ;
wire \ex_reg_rs2_bypass[16]~65_combout ;
wire \ex_reg_rs2_bypass[16]~66_combout ;
wire \alu_io_op2[16]~81_combout ;
wire \ex_reg_rs1_bypass[16]~66_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a16~portbdataout ;
wire \ex_rs_0~16_combout ;
wire \ex_rs_0[16]~q ;
wire \ex_reg_rs1_bypass[16]~67_combout ;
wire \ex_reg_rs1_bypass[16]~68_combout ;
wire \ex_reg_rs1_bypass[16]~69_combout ;
wire \alu_io_op1[16]~102_combout ;
wire \mem_alu_out~145_combout ;
wire \mem_alu_out~146_combout ;
wire \mem_alu_out~67_combout ;
wire \mem_alu_out~68_combout ;
wire \mem_alu_out~69_combout ;
wire \mem_alu_out[16]~q ;
wire \pc_cntr~52_combout ;
wire \pc_cntr~53_combout ;
wire \pc_cntr~54_combout ;
wire \pc_cntr[16]~q ;
wire \id_pc~15_combout ;
wire \ex_pc~15_combout ;
wire \ex_pc[17]~q ;
wire \npc[16]~29 ;
wire \npc[17]~30_combout ;
wire \id_npc~15_combout ;
wire \id_npc[17]~q ;
wire \ex_npc~15_combout ;
wire \ex_npc[17]~q ;
wire \mem_npc~13_combout ;
wire \mem_npc[17]~q ;
wire \wb_npc~13_combout ;
wire \wb_npc[17]~q ;
wire \mem_csr_data~22_combout ;
wire \mem_csr_data[17]~q ;
wire \wb_csr_data~15_combout ;
wire \wb_csr_data[17]~q ;
wire \wb_alu_out~15_combout ;
wire \wb_alu_out[17]~q ;
wire \_T_3543__T_3854_data[17]~33_combout ;
wire \wb_dmem_read_data~27_combout ;
wire \wb_dmem_read_data~29_combout ;
wire \wb_dmem_read_data~30_combout ;
wire \wb_dmem_read_data~76_combout ;
wire \wb_dmem_read_data[17]~q ;
wire \_T_3543__T_3854_data[17]~34_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a15~portbdataout ;
wire \ex_rs_0~17_combout ;
wire \ex_rs_0[17]~q ;
wire \ex_reg_rs1_bypass[17]~70_combout ;
wire \ex_reg_rs1_bypass[17]~71_combout ;
wire \ex_reg_rs1_bypass[17]~72_combout ;
wire \ex_reg_rs1_bypass[17]~73_combout ;
wire \alu_io_op1[17]~103_combout ;
wire \alu_io_op2[17]~56_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a15~portbdataout ;
wire \ex_rs_1~16_combout ;
wire \ex_rs_1[17]~q ;
wire \ex_reg_rs2_bypass[17]~59_combout ;
wire \ex_reg_rs2_bypass[17]~60_combout ;
wire \ex_reg_rs2_bypass[17]~61_combout ;
wire \ex_reg_rs2_bypass[17]~62_combout ;
wire \alu_io_op2[17]~80_combout ;
wire \mem_alu_out~70_combout ;
wire \mem_alu_out~71_combout ;
wire \mem_alu_out~72_combout ;
wire \mem_alu_out~73_combout ;
wire \mem_alu_out~74_combout ;
wire \mem_alu_out[17]~q ;
wire \mem_pc~15_combout ;
wire \mem_pc[17]~q ;
wire \mem_imm~32_combout ;
wire \mem_imm[17]~q ;
wire \_T_3862[16]~33 ;
wire \_T_3862[17]~34_combout ;
wire \pc_cntr~55_combout ;
wire \pc_cntr~56_combout ;
wire \pc_cntr~57_combout ;
wire \pc_cntr[17]~q ;
wire \id_pc~16_combout ;
wire \ex_pc~16_combout ;
wire \ex_pc[18]~q ;
wire \mem_pc~16_combout ;
wire \mem_pc[18]~q ;
wire \mem_imm~33_combout ;
wire \mem_imm[18]~q ;
wire \_T_3862[17]~35 ;
wire \_T_3862[18]~36_combout ;
wire \alu_io_op2[18]~58_combout ;
wire \mem_csr_data~23_combout ;
wire \mem_csr_data[18]~q ;
wire \wb_csr_data~16_combout ;
wire \wb_csr_data[18]~q ;
wire \npc[17]~31 ;
wire \npc[18]~32_combout ;
wire \id_npc~16_combout ;
wire \id_npc[18]~q ;
wire \ex_npc~16_combout ;
wire \ex_npc[18]~q ;
wire \mem_npc~14_combout ;
wire \mem_npc[18]~q ;
wire \wb_npc~14_combout ;
wire \wb_npc[18]~q ;
wire \wb_alu_out~16_combout ;
wire \wb_alu_out[18]~q ;
wire \_T_3543__T_3854_data[18]~35_combout ;
wire \wb_dmem_read_data~77_combout ;
wire \wb_dmem_read_data[18]~q ;
wire \_T_3543__T_3854_data[18]~36_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a14~portbdataout ;
wire \ex_rs_1~18_combout ;
wire \ex_rs_1[18]~q ;
wire \ex_reg_rs2_bypass[18]~67_combout ;
wire \ex_reg_rs2_bypass[18]~68_combout ;
wire \ex_reg_rs2_bypass[18]~69_combout ;
wire \ex_reg_rs2_bypass[18]~70_combout ;
wire \alu_io_op2[18]~82_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a14~portbdataout ;
wire \ex_rs_0~18_combout ;
wire \ex_rs_0[18]~q ;
wire \ex_reg_rs1_bypass[18]~74_combout ;
wire \ex_reg_rs1_bypass[18]~75_combout ;
wire \ex_reg_rs1_bypass[18]~76_combout ;
wire \ex_reg_rs1_bypass[18]~77_combout ;
wire \alu_io_op1[18]~104_combout ;
wire \mem_alu_out~75_combout ;
wire \mem_alu_out~76_combout ;
wire \mem_alu_out~77_combout ;
wire \mem_alu_out~78_combout ;
wire \mem_alu_out~79_combout ;
wire \mem_alu_out[18]~q ;
wire \pc_cntr~58_combout ;
wire \pc_cntr~59_combout ;
wire \pc_cntr~60_combout ;
wire \pc_cntr[18]~q ;
wire \id_pc~17_combout ;
wire \ex_pc~17_combout ;
wire \ex_pc[19]~q ;
wire \npc[18]~33 ;
wire \npc[19]~34_combout ;
wire \id_npc~17_combout ;
wire \id_npc[19]~q ;
wire \ex_npc~17_combout ;
wire \ex_npc[19]~q ;
wire \mem_npc~15_combout ;
wire \mem_npc[19]~q ;
wire \wb_npc~15_combout ;
wire \wb_npc[19]~q ;
wire \mem_csr_data~24_combout ;
wire \mem_csr_data[19]~q ;
wire \wb_csr_data~17_combout ;
wire \wb_csr_data[19]~q ;
wire \wb_alu_out~17_combout ;
wire \wb_alu_out[19]~q ;
wire \_T_3543__T_3854_data[19]~37_combout ;
wire \wb_dmem_read_data~78_combout ;
wire \wb_dmem_read_data[19]~q ;
wire \_T_3543__T_3854_data[19]~38_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a13~portbdataout ;
wire \ex_rs_0~19_combout ;
wire \ex_rs_0[19]~q ;
wire \ex_reg_rs1_bypass[19]~78_combout ;
wire \ex_reg_rs1_bypass[19]~79_combout ;
wire \ex_reg_rs1_bypass[19]~80_combout ;
wire \ex_reg_rs1_bypass[19]~81_combout ;
wire \alu_io_op1[19]~105_combout ;
wire \alu_io_op2[19]~59_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a13~portbdataout ;
wire \ex_rs_1~19_combout ;
wire \ex_rs_1[19]~q ;
wire \ex_reg_rs2_bypass[19]~71_combout ;
wire \ex_reg_rs2_bypass[19]~72_combout ;
wire \ex_reg_rs2_bypass[19]~73_combout ;
wire \ex_reg_rs2_bypass[19]~74_combout ;
wire \alu_io_op2[19]~93_combout ;
wire \mem_alu_out~80_combout ;
wire \mem_alu_out~81_combout ;
wire \mem_alu_out~82_combout ;
wire \mem_alu_out~83_combout ;
wire \mem_alu_out~84_combout ;
wire \mem_alu_out[19]~q ;
wire \mem_pc~17_combout ;
wire \mem_pc[19]~q ;
wire \mem_imm~34_combout ;
wire \mem_imm[19]~q ;
wire \_T_3862[18]~37 ;
wire \_T_3862[19]~38_combout ;
wire \pc_cntr~61_combout ;
wire \pc_cntr~62_combout ;
wire \pc_cntr~63_combout ;
wire \pc_cntr[19]~q ;
wire \id_pc~18_combout ;
wire \ex_pc~18_combout ;
wire \ex_pc[20]~q ;
wire \mem_pc~18_combout ;
wire \mem_pc[20]~q ;
wire \mem_imm~9_combout ;
wire \mem_imm~35_combout ;
wire \mem_imm[20]~q ;
wire \_T_3862[19]~39 ;
wire \_T_3862[20]~40_combout ;
wire \mem_csr_data~31_combout ;
wire \mem_csr_data[20]~q ;
wire \wb_csr_data~24_combout ;
wire \wb_csr_data[20]~q ;
wire \npc[19]~35 ;
wire \npc[20]~36_combout ;
wire \id_npc~24_combout ;
wire \id_npc[20]~q ;
wire \ex_npc~24_combout ;
wire \ex_npc[20]~q ;
wire \mem_npc~22_combout ;
wire \mem_npc[20]~q ;
wire \wb_npc~22_combout ;
wire \wb_npc[20]~q ;
wire \wb_alu_out~24_combout ;
wire \wb_alu_out[20]~q ;
wire \_T_3543__T_3854_data[20]~51_combout ;
wire \wb_dmem_read_data~79_combout ;
wire \wb_dmem_read_data[20]~q ;
wire \_T_3543__T_3854_data[20]~52_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a12~portbdataout ;
wire \ex_rs_1~27_combout ;
wire \ex_rs_1[20]~q ;
wire \ex_reg_rs2_bypass[20]~96_combout ;
wire \ex_reg_rs2_bypass[20]~97_combout ;
wire \ex_reg_rs2_bypass[20]~98_combout ;
wire \ex_reg_rs2_bypass[20]~99_combout ;
wire \alu_io_op2[20]~84_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a12~portbdataout ;
wire \ex_rs_0~26_combout ;
wire \ex_rs_0[20]~q ;
wire \ex_reg_rs1_bypass[20]~106_combout ;
wire \ex_reg_rs1_bypass[20]~107_combout ;
wire \ex_reg_rs1_bypass[20]~108_combout ;
wire \ex_reg_rs1_bypass[20]~109_combout ;
wire \alu_io_op1[20]~112_combout ;
wire \mem_alu_out~137_combout ;
wire \mem_alu_out~138_combout ;
wire \mem_alu_out~99_combout ;
wire \mem_alu_out~100_combout ;
wire \mem_alu_out~101_combout ;
wire \mem_alu_out[20]~q ;
wire \pc_cntr~64_combout ;
wire \pc_cntr~65_combout ;
wire \pc_cntr~66_combout ;
wire \pc_cntr[20]~q ;
wire \id_pc~19_combout ;
wire \ex_pc~19_combout ;
wire \ex_pc[21]~q ;
wire \npc[20]~37 ;
wire \npc[21]~38_combout ;
wire \id_npc~25_combout ;
wire \id_npc[21]~q ;
wire \ex_npc~25_combout ;
wire \ex_npc[21]~q ;
wire \mem_npc~23_combout ;
wire \mem_npc[21]~q ;
wire \wb_npc~23_combout ;
wire \wb_npc[21]~q ;
wire \mem_csr_data~37_combout ;
wire \mem_csr_data[21]~q ;
wire \wb_csr_data~25_combout ;
wire \wb_csr_data[21]~q ;
wire \wb_alu_out~25_combout ;
wire \wb_alu_out[21]~q ;
wire \_T_3543__T_3854_data[21]~53_combout ;
wire \wb_dmem_read_data~80_combout ;
wire \wb_dmem_read_data[21]~q ;
wire \_T_3543__T_3854_data[21]~54_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a11~portbdataout ;
wire \ex_rs_0~27_combout ;
wire \ex_rs_0[21]~q ;
wire \ex_reg_rs1_bypass[21]~110_combout ;
wire \ex_reg_rs1_bypass[21]~111_combout ;
wire \ex_reg_rs1_bypass[21]~112_combout ;
wire \ex_reg_rs1_bypass[21]~113_combout ;
wire \alu_io_op1[21]~113_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a11~portbdataout ;
wire \ex_rs_1~26_combout ;
wire \ex_rs_1[21]~q ;
wire \ex_reg_rs2_bypass[21]~92_combout ;
wire \ex_reg_rs2_bypass[21]~93_combout ;
wire \ex_reg_rs2_bypass[21]~94_combout ;
wire \ex_reg_rs2_bypass[21]~95_combout ;
wire \mem_imm~8_combout ;
wire \alu_io_op2[21]~83_combout ;
wire \mem_alu_out~102_combout ;
wire \mem_alu_out~103_combout ;
wire \mem_alu_out~104_combout ;
wire \mem_alu_out~105_combout ;
wire \mem_alu_out~106_combout ;
wire \mem_alu_out[21]~q ;
wire \mem_pc~19_combout ;
wire \mem_pc[21]~q ;
wire \mem_imm~36_combout ;
wire \mem_imm[21]~q ;
wire \_T_3862[20]~41 ;
wire \_T_3862[21]~42_combout ;
wire \pc_cntr~67_combout ;
wire \pc_cntr~68_combout ;
wire \pc_cntr~69_combout ;
wire \pc_cntr[21]~q ;
wire \id_pc~20_combout ;
wire \ex_pc~20_combout ;
wire \ex_pc[22]~q ;
wire \mem_pc~20_combout ;
wire \mem_pc[22]~q ;
wire \mem_imm~10_combout ;
wire \mem_imm~37_combout ;
wire \mem_imm[22]~q ;
wire \_T_3862[21]~43 ;
wire \_T_3862[22]~44_combout ;
wire \mem_csr_data~32_combout ;
wire \mem_csr_data[22]~q ;
wire \wb_csr_data~26_combout ;
wire \wb_csr_data[22]~q ;
wire \npc[21]~39 ;
wire \npc[22]~40_combout ;
wire \id_npc~26_combout ;
wire \id_npc[22]~q ;
wire \ex_npc~26_combout ;
wire \ex_npc[22]~q ;
wire \mem_npc~24_combout ;
wire \mem_npc[22]~q ;
wire \wb_npc~24_combout ;
wire \wb_npc[22]~q ;
wire \wb_alu_out~26_combout ;
wire \wb_alu_out[22]~q ;
wire \_T_3543__T_3854_data[22]~55_combout ;
wire \wb_dmem_read_data~81_combout ;
wire \wb_dmem_read_data[22]~q ;
wire \_T_3543__T_3854_data[22]~56_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a10~portbdataout ;
wire \ex_rs_1~28_combout ;
wire \ex_rs_1[22]~q ;
wire \ex_reg_rs2_bypass[22]~100_combout ;
wire \ex_reg_rs2_bypass[22]~101_combout ;
wire \ex_reg_rs2_bypass[22]~102_combout ;
wire \ex_reg_rs2_bypass[22]~103_combout ;
wire \alu_io_op2[22]~85_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a10~portbdataout ;
wire \ex_rs_0~28_combout ;
wire \ex_rs_0[22]~q ;
wire \ex_reg_rs1_bypass[22]~114_combout ;
wire \ex_reg_rs1_bypass[22]~115_combout ;
wire \ex_reg_rs1_bypass[22]~116_combout ;
wire \ex_reg_rs1_bypass[22]~117_combout ;
wire \alu_io_op1[22]~114_combout ;
wire \mem_alu_out~135_combout ;
wire \mem_alu_out~136_combout ;
wire \mem_alu_out~107_combout ;
wire \mem_alu_out~108_combout ;
wire \mem_alu_out~109_combout ;
wire \mem_alu_out[22]~q ;
wire \pc_cntr~70_combout ;
wire \pc_cntr~71_combout ;
wire \pc_cntr~72_combout ;
wire \pc_cntr[22]~q ;
wire \id_pc~21_combout ;
wire \ex_pc~21_combout ;
wire \ex_pc[23]~q ;
wire \npc[22]~41 ;
wire \npc[23]~42_combout ;
wire \id_npc~27_combout ;
wire \id_npc[23]~q ;
wire \ex_npc~27_combout ;
wire \ex_npc[23]~q ;
wire \mem_npc~25_combout ;
wire \mem_npc[23]~q ;
wire \wb_npc~25_combout ;
wire \wb_npc[23]~q ;
wire \mem_csr_data~33_combout ;
wire \mem_csr_data[23]~q ;
wire \wb_csr_data~27_combout ;
wire \wb_csr_data[23]~q ;
wire \wb_alu_out~27_combout ;
wire \wb_alu_out[23]~q ;
wire \_T_3543__T_3854_data[23]~57_combout ;
wire \wb_dmem_read_data~82_combout ;
wire \wb_dmem_read_data~83_combout ;
wire \wb_dmem_read_data~84_combout ;
wire \wb_dmem_read_data[23]~q ;
wire \_T_3543__T_3854_data[23]~58_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a9~portbdataout ;
wire \ex_rs_0~29_combout ;
wire \ex_rs_0[23]~q ;
wire \ex_reg_rs1_bypass[23]~118_combout ;
wire \ex_reg_rs1_bypass[23]~119_combout ;
wire \ex_reg_rs1_bypass[23]~120_combout ;
wire \ex_reg_rs1_bypass[23]~121_combout ;
wire \alu_io_op1[23]~119_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a9~portbdataout ;
wire \ex_rs_1~29_combout ;
wire \ex_rs_1[23]~q ;
wire \ex_reg_rs2_bypass[23]~104_combout ;
wire \ex_reg_rs2_bypass[23]~105_combout ;
wire \ex_reg_rs2_bypass[23]~106_combout ;
wire \ex_reg_rs2_bypass[23]~107_combout ;
wire \mem_imm~11_combout ;
wire \alu_io_op2[23]~86_combout ;
wire \mem_alu_out~110_combout ;
wire \mem_alu_out~111_combout ;
wire \mem_alu_out~112_combout ;
wire \mem_alu_out~113_combout ;
wire \mem_alu_out~114_combout ;
wire \mem_alu_out[23]~q ;
wire \mem_pc~21_combout ;
wire \mem_pc[23]~q ;
wire \mem_imm~38_combout ;
wire \mem_imm[23]~q ;
wire \_T_3862[22]~45 ;
wire \_T_3862[23]~46_combout ;
wire \pc_cntr~73_combout ;
wire \pc_cntr~74_combout ;
wire \pc_cntr~75_combout ;
wire \pc_cntr[23]~q ;
wire \id_pc~22_combout ;
wire \ex_pc~22_combout ;
wire \ex_pc[24]~q ;
wire \mem_pc~22_combout ;
wire \mem_pc[24]~q ;
wire \mem_imm~13_combout ;
wire \mem_imm~39_combout ;
wire \mem_imm[24]~q ;
wire \_T_3862[23]~47 ;
wire \_T_3862[24]~48_combout ;
wire \mem_csr_data~34_combout ;
wire \mem_csr_data[24]~q ;
wire \wb_csr_data~28_combout ;
wire \wb_csr_data[24]~q ;
wire \npc[23]~43 ;
wire \npc[24]~44_combout ;
wire \id_npc~28_combout ;
wire \id_npc[24]~q ;
wire \ex_npc~28_combout ;
wire \ex_npc[24]~q ;
wire \mem_npc~26_combout ;
wire \mem_npc[24]~q ;
wire \wb_npc~26_combout ;
wire \wb_npc[24]~q ;
wire \wb_alu_out~28_combout ;
wire \wb_alu_out[24]~q ;
wire \_T_3543__T_3854_data[24]~59_combout ;
wire \wb_dmem_read_data~85_combout ;
wire \wb_dmem_read_data[24]~q ;
wire \_T_3543__T_3854_data[24]~60_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a8~portbdataout ;
wire \ex_rs_1~31_combout ;
wire \ex_rs_1[24]~q ;
wire \ex_reg_rs2_bypass[24]~112_combout ;
wire \ex_reg_rs2_bypass[24]~113_combout ;
wire \ex_reg_rs2_bypass[24]~114_combout ;
wire \ex_reg_rs2_bypass[24]~115_combout ;
wire \alu_io_op2[24]~88_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a8~portbdataout ;
wire \ex_rs_0~30_combout ;
wire \ex_rs_0[24]~q ;
wire \ex_reg_rs1_bypass[24]~122_combout ;
wire \ex_reg_rs1_bypass[24]~123_combout ;
wire \ex_reg_rs1_bypass[24]~124_combout ;
wire \ex_reg_rs1_bypass[24]~125_combout ;
wire \alu_io_op1[24]~115_combout ;
wire \mem_alu_out~133_combout ;
wire \mem_alu_out~134_combout ;
wire \mem_alu_out~115_combout ;
wire \mem_alu_out~116_combout ;
wire \mem_alu_out~117_combout ;
wire \mem_alu_out[24]~q ;
wire \pc_cntr~76_combout ;
wire \pc_cntr~77_combout ;
wire \pc_cntr~78_combout ;
wire \pc_cntr[24]~q ;
wire \id_pc~23_combout ;
wire \ex_pc~23_combout ;
wire \ex_pc[25]~q ;
wire \npc[24]~45 ;
wire \npc[25]~46_combout ;
wire \id_npc~29_combout ;
wire \id_npc[25]~q ;
wire \ex_npc~29_combout ;
wire \ex_npc[25]~q ;
wire \mem_npc~27_combout ;
wire \mem_npc[25]~q ;
wire \wb_npc~27_combout ;
wire \wb_npc[25]~q ;
wire \mem_csr_data~38_combout ;
wire \mem_csr_data[25]~q ;
wire \wb_csr_data~29_combout ;
wire \wb_csr_data[25]~q ;
wire \wb_alu_out~29_combout ;
wire \wb_alu_out[25]~q ;
wire \_T_3543__T_3854_data[25]~61_combout ;
wire \wb_dmem_read_data~86_combout ;
wire \wb_dmem_read_data[25]~q ;
wire \_T_3543__T_3854_data[25]~62_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a7~portbdataout ;
wire \ex_rs_0~31_combout ;
wire \ex_rs_0[25]~q ;
wire \ex_reg_rs1_bypass[25]~126_combout ;
wire \ex_reg_rs1_bypass[25]~127_combout ;
wire \ex_reg_rs1_bypass[25]~128_combout ;
wire \ex_reg_rs1_bypass[25]~129_combout ;
wire \alu_io_op1[25]~116_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a7~portbdataout ;
wire \ex_rs_1~30_combout ;
wire \ex_rs_1[25]~q ;
wire \ex_reg_rs2_bypass[25]~108_combout ;
wire \ex_reg_rs2_bypass[25]~109_combout ;
wire \ex_reg_rs2_bypass[25]~110_combout ;
wire \ex_reg_rs2_bypass[25]~111_combout ;
wire \mem_imm~12_combout ;
wire \alu_io_op2[25]~87_combout ;
wire \mem_alu_out~118_combout ;
wire \mem_alu_out~119_combout ;
wire \mem_alu_out~120_combout ;
wire \mem_alu_out~121_combout ;
wire \mem_alu_out~122_combout ;
wire \mem_alu_out[25]~q ;
wire \mem_pc~23_combout ;
wire \mem_pc[25]~q ;
wire \mem_imm~40_combout ;
wire \mem_imm[25]~q ;
wire \_T_3862[24]~49 ;
wire \_T_3862[25]~50_combout ;
wire \pc_cntr~79_combout ;
wire \pc_cntr~80_combout ;
wire \pc_cntr~81_combout ;
wire \pc_cntr[25]~q ;
wire \id_pc~24_combout ;
wire \ex_pc~24_combout ;
wire \ex_pc[26]~q ;
wire \mem_pc~24_combout ;
wire \mem_pc[26]~q ;
wire \mem_imm~14_combout ;
wire \mem_imm~41_combout ;
wire \mem_imm[26]~q ;
wire \_T_3862[25]~51 ;
wire \_T_3862[26]~52_combout ;
wire \mem_csr_data~35_combout ;
wire \mem_csr_data[26]~q ;
wire \wb_csr_data~30_combout ;
wire \wb_csr_data[26]~q ;
wire \npc[25]~47 ;
wire \npc[26]~48_combout ;
wire \id_npc~30_combout ;
wire \id_npc[26]~q ;
wire \ex_npc~30_combout ;
wire \ex_npc[26]~q ;
wire \mem_npc~28_combout ;
wire \mem_npc[26]~q ;
wire \wb_npc~28_combout ;
wire \wb_npc[26]~q ;
wire \wb_alu_out~30_combout ;
wire \wb_alu_out[26]~q ;
wire \_T_3543__T_3854_data[26]~63_combout ;
wire \wb_dmem_read_data~87_combout ;
wire \wb_dmem_read_data[26]~q ;
wire \_T_3543__T_3854_data[26]~64_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a6~portbdataout ;
wire \ex_rs_1~32_combout ;
wire \ex_rs_1[26]~q ;
wire \ex_reg_rs2_bypass[26]~116_combout ;
wire \ex_reg_rs2_bypass[26]~117_combout ;
wire \ex_reg_rs2_bypass[26]~118_combout ;
wire \ex_reg_rs2_bypass[26]~119_combout ;
wire \alu_io_op2[26]~89_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a6~portbdataout ;
wire \ex_rs_0~32_combout ;
wire \ex_rs_0[26]~q ;
wire \ex_reg_rs1_bypass[26]~130_combout ;
wire \ex_reg_rs1_bypass[26]~131_combout ;
wire \ex_reg_rs1_bypass[26]~132_combout ;
wire \ex_reg_rs1_bypass[26]~133_combout ;
wire \alu_io_op1[26]~117_combout ;
wire \mem_alu_out~131_combout ;
wire \mem_alu_out~132_combout ;
wire \mem_alu_out~123_combout ;
wire \mem_alu_out~124_combout ;
wire \mem_alu_out~125_combout ;
wire \mem_alu_out[26]~q ;
wire \pc_cntr~82_combout ;
wire \pc_cntr~83_combout ;
wire \pc_cntr~84_combout ;
wire \pc_cntr[26]~q ;
wire \id_pc~25_combout ;
wire \ex_pc~25_combout ;
wire \ex_pc[27]~q ;
wire \npc[26]~49 ;
wire \npc[27]~50_combout ;
wire \id_npc~31_combout ;
wire \id_npc[27]~q ;
wire \ex_npc~31_combout ;
wire \ex_npc[27]~q ;
wire \mem_npc~29_combout ;
wire \mem_npc[27]~q ;
wire \wb_npc~29_combout ;
wire \wb_npc[27]~q ;
wire \mem_csr_data~39_combout ;
wire \mem_csr_data[27]~q ;
wire \wb_csr_data~31_combout ;
wire \wb_csr_data[27]~q ;
wire \wb_alu_out~31_combout ;
wire \wb_alu_out[27]~q ;
wire \_T_3543__T_3854_data[27]~65_combout ;
wire \wb_dmem_read_data~88_combout ;
wire \wb_dmem_read_data[27]~q ;
wire \_T_3543__T_3854_data[27]~66_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a5~portbdataout ;
wire \ex_rs_0~33_combout ;
wire \ex_rs_0[27]~q ;
wire \ex_reg_rs1_bypass[27]~134_combout ;
wire \ex_reg_rs1_bypass[27]~135_combout ;
wire \ex_reg_rs1_bypass[27]~136_combout ;
wire \ex_reg_rs1_bypass[27]~137_combout ;
wire \alu_io_op1[27]~118_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a5~portbdataout ;
wire \ex_rs_1~33_combout ;
wire \ex_rs_1[27]~q ;
wire \ex_reg_rs2_bypass[27]~120_combout ;
wire \ex_reg_rs2_bypass[27]~121_combout ;
wire \ex_reg_rs2_bypass[27]~122_combout ;
wire \ex_reg_rs2_bypass[27]~123_combout ;
wire \mem_imm~15_combout ;
wire \alu_io_op2[27]~90_combout ;
wire \mem_alu_out~126_combout ;
wire \mem_alu_out~127_combout ;
wire \mem_alu_out~128_combout ;
wire \mem_alu_out~129_combout ;
wire \mem_alu_out~130_combout ;
wire \mem_alu_out[27]~q ;
wire \mem_pc~25_combout ;
wire \mem_pc[27]~q ;
wire \mem_imm~42_combout ;
wire \mem_imm[27]~q ;
wire \_T_3862[26]~53 ;
wire \_T_3862[27]~54_combout ;
wire \pc_cntr~85_combout ;
wire \pc_cntr~86_combout ;
wire \pc_cntr~87_combout ;
wire \pc_cntr[27]~q ;
wire \id_pc~26_combout ;
wire \ex_pc~26_combout ;
wire \ex_pc[28]~q ;
wire \mem_pc~26_combout ;
wire \mem_pc[28]~q ;
wire \mem_imm~5_combout ;
wire \mem_imm~43_combout ;
wire \mem_imm[28]~q ;
wire \_T_3862[27]~55 ;
wire \_T_3862[28]~56_combout ;
wire \mem_csr_data~10_combout ;
wire \mem_csr_data[28]~q ;
wire \wb_csr_data~2_combout ;
wire \wb_csr_data[28]~q ;
wire \npc[27]~51 ;
wire \npc[28]~52_combout ;
wire \id_npc~2_combout ;
wire \id_npc[28]~q ;
wire \ex_npc~2_combout ;
wire \ex_npc[28]~q ;
wire \mem_npc~0_combout ;
wire \mem_npc[28]~q ;
wire \wb_npc~0_combout ;
wire \wb_npc[28]~q ;
wire \wb_alu_out~2_combout ;
wire \wb_alu_out[28]~q ;
wire \_T_3543__T_3854_data[28]~7_combout ;
wire \wb_dmem_read_data~33_combout ;
wire \wb_dmem_read_data[28]~q ;
wire \_T_3543__T_3854_data[28]~8_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a4~portbdataout ;
wire \ex_rs_1~5_combout ;
wire \ex_rs_1[28]~q ;
wire \ex_reg_rs2_bypass[28]~19_combout ;
wire \ex_reg_rs2_bypass[28]~20_combout ;
wire \ex_reg_rs2_bypass[28]~21_combout ;
wire \ex_reg_rs2_bypass[28]~22_combout ;
wire \alu_io_op2[28]~74_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a4~portbdataout ;
wire \ex_rs_0~4_combout ;
wire \ex_rs_0[28]~q ;
wire \ex_reg_rs1_bypass[28]~17_combout ;
wire \ex_reg_rs1_bypass[28]~18_combout ;
wire \ex_reg_rs1_bypass[28]~19_combout ;
wire \ex_reg_rs1_bypass[28]~21_combout ;
wire \alu_io_op1[28]~90_combout ;
wire \mem_alu_out~159_combout ;
wire \mem_alu_out~160_combout ;
wire \mem_alu_out~21_combout ;
wire \mem_alu_out~22_combout ;
wire \mem_alu_out~23_combout ;
wire \mem_alu_out[28]~q ;
wire \pc_cntr~88_combout ;
wire \pc_cntr~89_combout ;
wire \pc_cntr~90_combout ;
wire \pc_cntr[28]~q ;
wire \id_pc~27_combout ;
wire \ex_pc~27_combout ;
wire \ex_pc[29]~q ;
wire \npc[28]~53 ;
wire \npc[29]~54_combout ;
wire \id_npc~3_combout ;
wire \id_npc[29]~q ;
wire \ex_npc~3_combout ;
wire \ex_npc[29]~q ;
wire \mem_npc~1_combout ;
wire \mem_npc[29]~q ;
wire \wb_npc~1_combout ;
wire \wb_npc[29]~q ;
wire \mem_csr_data~36_combout ;
wire \mem_csr_data[29]~q ;
wire \wb_csr_data~3_combout ;
wire \wb_csr_data[29]~q ;
wire \wb_alu_out~3_combout ;
wire \wb_alu_out[29]~q ;
wire \_T_3543__T_3854_data[29]~9_combout ;
wire \wb_dmem_read_data~37_combout ;
wire \wb_dmem_read_data[29]~q ;
wire \_T_3543__T_3854_data[29]~10_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a3~portbdataout ;
wire \ex_rs_0~5_combout ;
wire \ex_rs_0[29]~q ;
wire \ex_reg_rs1_bypass[29]~22_combout ;
wire \ex_reg_rs1_bypass[29]~23_combout ;
wire \ex_reg_rs1_bypass[29]~24_combout ;
wire \ex_reg_rs1_bypass[29]~25_combout ;
wire \alu_io_op1[29]~91_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a3~portbdataout ;
wire \ex_rs_1~4_combout ;
wire \ex_rs_1[29]~q ;
wire \ex_reg_rs2_bypass[29]~15_combout ;
wire \ex_reg_rs2_bypass[29]~16_combout ;
wire \ex_reg_rs2_bypass[29]~17_combout ;
wire \ex_reg_rs2_bypass[29]~18_combout ;
wire \mem_imm~4_combout ;
wire \alu_io_op2[29]~73_combout ;
wire \mem_alu_out~24_combout ;
wire \mem_alu_out~25_combout ;
wire \mem_alu_out~26_combout ;
wire \mem_alu_out~27_combout ;
wire \mem_alu_out~28_combout ;
wire \mem_alu_out[29]~q ;
wire \mem_pc~27_combout ;
wire \mem_pc[29]~q ;
wire \mem_imm~44_combout ;
wire \mem_imm[29]~q ;
wire \_T_3862[28]~57 ;
wire \_T_3862[29]~58_combout ;
wire \pc_cntr~91_combout ;
wire \pc_cntr~92_combout ;
wire \pc_cntr~93_combout ;
wire \pc_cntr[29]~q ;
wire \id_pc~28_combout ;
wire \ex_pc~28_combout ;
wire \ex_pc[30]~q ;
wire \mem_pc~28_combout ;
wire \mem_pc[30]~q ;
wire \mem_imm~6_combout ;
wire \mem_imm~45_combout ;
wire \mem_imm[30]~q ;
wire \_T_3862[29]~59 ;
wire \_T_3862[30]~60_combout ;
wire \mem_csr_data~11_combout ;
wire \mem_csr_data[30]~q ;
wire \wb_csr_data~4_combout ;
wire \wb_csr_data[30]~q ;
wire \npc[29]~55 ;
wire \npc[30]~56_combout ;
wire \id_npc~4_combout ;
wire \id_npc[30]~q ;
wire \ex_npc~4_combout ;
wire \ex_npc[30]~q ;
wire \mem_npc~2_combout ;
wire \mem_npc[30]~q ;
wire \wb_npc~2_combout ;
wire \wb_npc[30]~q ;
wire \wb_alu_out~4_combout ;
wire \wb_alu_out[30]~q ;
wire \_T_3543__T_3854_data[30]~11_combout ;
wire \wb_dmem_read_data~38_combout ;
wire \wb_dmem_read_data[30]~q ;
wire \_T_3543__T_3854_data[30]~12_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a2~portbdataout ;
wire \ex_rs_1~6_combout ;
wire \ex_rs_1[30]~q ;
wire \ex_reg_rs2_bypass[30]~23_combout ;
wire \ex_reg_rs2_bypass[30]~24_combout ;
wire \ex_reg_rs2_bypass[30]~25_combout ;
wire \ex_reg_rs2_bypass[30]~26_combout ;
wire \alu_io_op2[30]~75_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a2~portbdataout ;
wire \ex_rs_0~6_combout ;
wire \ex_rs_0[30]~q ;
wire \ex_reg_rs1_bypass[30]~26_combout ;
wire \ex_reg_rs1_bypass[30]~27_combout ;
wire \ex_reg_rs1_bypass[30]~28_combout ;
wire \ex_reg_rs1_bypass[30]~29_combout ;
wire \alu_io_op1[30]~92_combout ;
wire \mem_alu_out~157_combout ;
wire \mem_alu_out~158_combout ;
wire \mem_alu_out~29_combout ;
wire \mem_alu_out~30_combout ;
wire \mem_alu_out~31_combout ;
wire \mem_alu_out[30]~q ;
wire \pc_cntr~94_combout ;
wire \pc_cntr~95_combout ;
wire \pc_cntr~96_combout ;
wire \pc_cntr[30]~q ;
wire \id_pc~29_combout ;
wire \ex_pc~29_combout ;
wire \ex_pc[31]~q ;
wire \npc[30]~57 ;
wire \npc[31]~58_combout ;
wire \id_npc~5_combout ;
wire \id_npc[31]~q ;
wire \ex_npc~5_combout ;
wire \ex_npc[31]~q ;
wire \mem_npc~3_combout ;
wire \mem_npc[31]~q ;
wire \wb_npc~3_combout ;
wire \wb_npc[31]~q ;
wire \mem_csr_data~12_combout ;
wire \mem_csr_data[31]~q ;
wire \wb_csr_data~5_combout ;
wire \wb_csr_data[31]~q ;
wire \wb_alu_out~5_combout ;
wire \wb_alu_out[31]~q ;
wire \_T_3543__T_3854_data[31]~13_combout ;
wire \wb_dmem_read_data~40_combout ;
wire \wb_dmem_read_data~41_combout ;
wire \wb_dmem_read_data~42_combout ;
wire \wb_dmem_read_data[31]~q ;
wire \_T_3543__T_3854_data[31]~14_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a1~portbdataout ;
wire \ex_rs_0~7_combout ;
wire \ex_rs_0[31]~q ;
wire \ex_reg_rs1_bypass[31]~30_combout ;
wire \ex_reg_rs1_bypass[31]~31_combout ;
wire \ex_reg_rs1_bypass[31]~32_combout ;
wire \ex_reg_rs1_bypass[31]~33_combout ;
wire \alu_io_op1[31]~93_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a1~portbdataout ;
wire \ex_rs_1~7_combout ;
wire \ex_rs_1[31]~q ;
wire \ex_reg_rs2_bypass[31]~27_combout ;
wire \ex_reg_rs2_bypass[31]~28_combout ;
wire \ex_reg_rs2_bypass[31]~29_combout ;
wire \ex_reg_rs2_bypass[31]~30_combout ;
wire \alu_io_op2[31]~76_combout ;
wire \mem_alu_out~32_combout ;
wire \mem_alu_out~33_combout ;
wire \mem_alu_out~34_combout ;
wire \mem_alu_out~35_combout ;
wire \mem_alu_out~36_combout ;
wire \mem_alu_out[31]~q ;
wire \mem_pc~29_combout ;
wire \mem_pc[31]~q ;
wire \mem_imm~47_combout ;
wire \mem_imm[31]~q ;
wire \_T_3862[30]~61 ;
wire \_T_3862[31]~62_combout ;
wire \pc_cntr~97_combout ;
wire \pc_cntr~98_combout ;
wire \pc_cntr~99_combout ;
wire \pc_cntr[31]~q ;
wire \id_pc~30_combout ;
wire \mem_csr_data~8_combout ;
wire \mem_csr_data[1]~q ;
wire \ex_reg_rs2_bypass[1]~126_combout ;
wire \wb_alu_out~0_combout ;
wire \wb_alu_out[1]~q ;
wire \wb_csr_data~0_combout ;
wire \wb_csr_data[1]~q ;
wire \_T_3543__T_3854_data[23]~0_combout ;
wire \wb_dmem_read_data[1]~7_combout ;
wire \wb_dmem_read_data[1]~q ;
wire \_T_3543__T_3854_data[1]~3_combout ;
wire \_T_3543__T_3854_data[1]~4_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a31~portbdataout ;
wire \ex_rs_1~2_combout ;
wire \ex_rs_1[1]~q ;
wire \ex_reg_rs2_bypass[1]~6_combout ;
wire \ex_reg_rs2_bypass[1]~7_combout ;
wire \ex_reg_rs2_bypass[1]~8_combout ;
wire \ex_reg_rs2_bypass[1]~9_combout ;
wire \csr_io_alu_op2[1]~1_combout ;
wire \_T_3639~0_combout ;
wire \ex_reg_rs1_bypass[1]~5_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a31~portbdataout ;
wire \ex_rs_0~2_combout ;
wire \ex_rs_0[1]~q ;
wire \ex_reg_rs1_bypass[1]~9_combout ;
wire \ex_reg_rs1_bypass[1]~10_combout ;
wire \ex_reg_rs1_bypass[1]~11_combout ;
wire \ex_npc~1_combout ;
wire \ex_npc[1]~q ;
wire \csr_io_alu_op1[1]~7_combout ;
wire \mem_alu_out~163_combout ;
wire \mem_alu_out~164_combout ;
wire \mem_alu_out~3_combout ;
wire \mem_alu_out~4_combout ;
wire \mem_alu_out~7_combout ;
wire \mem_csr_data~9_combout ;
wire \mem_csr_data[0]~q ;
wire \ex_reg_rs1_bypass[0]~13_combout ;
wire \wb_csr_data~1_combout ;
wire \wb_csr_data[0]~q ;
wire \wb_alu_out~1_combout ;
wire \wb_alu_out[0]~q ;
wire \_T_3543__T_3854_data[0]~5_combout ;
wire \wb_dmem_read_data[0]~0_combout ;
wire \wb_dmem_read_data[0]~q ;
wire \_T_3543__T_3854_data[0]~6_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a0~portbdataout ;
wire \ex_rs_0~3_combout ;
wire \ex_rs_0[0]~q ;
wire \ex_reg_rs1_bypass[0]~14_combout ;
wire \ex_reg_rs1_bypass[0]~15_combout ;
wire \ex_reg_rs1_bypass[0]~16_combout ;
wire \ex_npc~0_combout ;
wire \ex_npc[0]~q ;
wire \csr_io_alu_op1[0]~8_combout ;
wire \mem_alu_out~8_combout ;
wire \mem_alu_out~9_combout ;
wire \csr_io_alu_op2[0]~2_combout ;
wire \alu_io_op2[3]~42_combout ;
wire \ex_reg_rs2_bypass[0]~10_combout ;
wire \ex_reg_rs2_bypass[0]~11_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a0~portbdataout ;
wire \ex_rs_1~3_combout ;
wire \ex_rs_1[0]~q ;
wire \ex_reg_rs2_bypass[0]~12_combout ;
wire \ex_reg_rs2_bypass[0]~13_combout ;
wire \ex_reg_rs2_bypass[0]~14_combout ;
wire \csr_io_alu_op2[0]~3_combout ;
wire \mem_alu_out~10_combout ;
wire \mem_alu_out~11_combout ;
wire \mem_alu_out~12_combout ;
wire \mem_ctrl_mem_wr~8_combout ;
wire \mem_rs_1~42_combout ;
wire \mem_csr_data~26_combout ;
wire \mem_csr_data[2]~q ;
wire \ex_reg_rs1_bypass[2]~86_combout ;
wire \wb_csr_data~19_combout ;
wire \wb_csr_data[2]~q ;
wire \id_npc~19_combout ;
wire \id_npc[2]~q ;
wire \ex_npc~19_combout ;
wire \ex_npc[2]~q ;
wire \mem_npc~17_combout ;
wire \mem_npc[2]~q ;
wire \wb_npc~17_combout ;
wire \wb_npc[2]~q ;
wire \wb_alu_out~19_combout ;
wire \wb_alu_out[2]~q ;
wire \_T_3543__T_3854_data[2]~41_combout ;
wire \wb_dmem_read_data[2]~6_combout ;
wire \wb_dmem_read_data[2]~q ;
wire \_T_3543__T_3854_data[2]~42_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a30~portbdataout ;
wire \ex_rs_0~21_combout ;
wire \ex_rs_0[2]~q ;
wire \ex_reg_rs1_bypass[2]~87_combout ;
wire \ex_reg_rs1_bypass[2]~88_combout ;
wire \ex_reg_rs1_bypass[2]~89_combout ;
wire \alu_io_op1[2]~107_combout ;
wire \ex_reg_rs2_bypass[2]~77_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a30~portbdataout ;
wire \ex_rs_1~21_combout ;
wire \ex_rs_1[2]~q ;
wire \ex_reg_rs2_bypass[2]~78_combout ;
wire \ex_reg_rs2_bypass[2]~79_combout ;
wire \ex_reg_rs2_bypass[2]~80_combout ;
wire \alu_io_op2[2]~63_combout ;
wire \alu_io_op2[2]~91_combout ;
wire \mem_alu_out~13_combout ;
wire \mem_alu_out~14_combout ;
wire \mem_alu_out~15_combout ;
wire \mem_alu_out~16_combout ;
wire \mem_alu_out~17_combout ;
wire \mem_csr_data~27_combout ;
wire \mem_csr_data[3]~q ;
wire \wb_alu_out~20_combout ;
wire \wb_alu_out[3]~q ;
wire \wb_csr_data~20_combout ;
wire \wb_csr_data[3]~q ;
wire \id_npc~20_combout ;
wire \id_npc[3]~q ;
wire \ex_npc~20_combout ;
wire \ex_npc[3]~q ;
wire \mem_npc~18_combout ;
wire \mem_npc[3]~q ;
wire \wb_npc~18_combout ;
wire \wb_npc[3]~q ;
wire \_T_3543__T_3854_data[3]~43_combout ;
wire \wb_dmem_read_data[3]~5_combout ;
wire \wb_dmem_read_data[3]~q ;
wire \_T_3543__T_3854_data[3]~44_combout ;
wire \_T_3543_rtl_0|auto_generated|ram_block1a29~portbdataout ;
wire \ex_rs_1~22_combout ;
wire \ex_rs_1[3]~q ;
wire \ex_reg_rs2_bypass[3]~81_combout ;
wire \ex_reg_rs2_bypass[3]~82_combout ;
wire \alu_io_op2[3]~64_combout ;
wire \alu_io_op2[3]~65_combout ;
wire \alu_io_op2[3]~66_combout ;
wire \ex_reg_rs1_bypass[3]~94_combout ;
wire \_T_3543_rtl_1|auto_generated|ram_block1a29~portbdataout ;
wire \ex_rs_0~23_combout ;
wire \ex_rs_0[3]~q ;
wire \ex_reg_rs1_bypass[3]~95_combout ;
wire \ex_reg_rs1_bypass[3]~96_combout ;
wire \ex_reg_rs1_bypass[3]~97_combout ;
wire \alu_io_op1[3]~109_combout ;
wire \mem_alu_out~161_combout ;
wire \mem_alu_out~162_combout ;
wire \mem_alu_out~18_combout ;
wire \mem_alu_out~19_combout ;
wire \mem_alu_out~20_combout ;
wire \mem_rs_1~43_combout ;
wire \mem_rs_1~53_combout ;
wire \ex_reg_rs2_bypass[3]~124_combout ;
wire \mem_rs_1~44_combout ;
wire \ex_reg_rs2_bypass[4]~125_combout ;
wire \mem_rs_1~45_combout ;
wire \mem_rs_1~46_combout ;
wire \mem_rs_1~47_combout ;
wire \mem_rs_1~48_combout ;
wire \mem_rs_1~49_combout ;
wire \mem_rs_1~50_combout ;
wire \mem_rs_1~51_combout ;
wire \mem_rs_1~52_combout ;
wire \mem_rs_1~54_combout ;
wire \mem_rs_1~55_combout ;
wire \mem_rs_1~56_combout ;
wire \mem_rs_1~57_combout ;
wire \mem_rs_1~58_combout ;
wire \mem_rs_1~59_combout ;
wire \mem_rs_1~60_combout ;
wire \mem_rs_1~61_combout ;
wire \mem_rs_1~62_combout ;
wire \mem_rs_1~63_combout ;
wire \mem_rs_1~64_combout ;
wire \mem_rs_1~65_combout ;
wire \ex_ctrl_mem_wr~12_combout ;
wire \ex_ctrl_mem_wr.00~q ;
wire \mem_ctrl_mem_wr~9_combout ;
wire \w_req~0_combout ;
wire \ex_ctrl_mem_wr~11_combout ;
wire \ex_ctrl_mem_wr~13_combout ;
wire \ex_ctrl_mem_wr.01~q ;
wire \mem_ctrl_mem_wr~10_combout ;
wire \io_w_dmem_dat_data[24]~32_combout ;
wire \mem_rs_1~66_combout ;
wire \mem_rs_1[24]~q ;
wire \io_w_dmem_dat_data[24]~33_combout ;
wire \io_w_dmem_dat_data[25]~34_combout ;
wire \mem_rs_1~67_combout ;
wire \mem_rs_1[25]~q ;
wire \io_w_dmem_dat_data[25]~35_combout ;
wire \io_w_dmem_dat_data[26]~36_combout ;
wire \mem_rs_1~68_combout ;
wire \mem_rs_1[26]~q ;
wire \io_w_dmem_dat_data[26]~37_combout ;
wire \io_w_dmem_dat_data[27]~38_combout ;
wire \mem_rs_1~69_combout ;
wire \mem_rs_1[27]~q ;
wire \io_w_dmem_dat_data[27]~39_combout ;
wire \io_w_dmem_dat_data[28]~40_combout ;
wire \mem_rs_1~70_combout ;
wire \mem_rs_1[28]~q ;
wire \io_w_dmem_dat_data[28]~41_combout ;
wire \io_w_dmem_dat_data[29]~42_combout ;
wire \mem_rs_1~71_combout ;
wire \mem_rs_1[29]~q ;
wire \io_w_dmem_dat_data[29]~43_combout ;
wire \io_w_dmem_dat_data[30]~44_combout ;
wire \mem_rs_1~72_combout ;
wire \mem_rs_1[30]~q ;
wire \io_w_dmem_dat_data[30]~45_combout ;
wire \io_w_dmem_dat_data[31]~46_combout ;
wire \mem_rs_1~73_combout ;
wire \mem_rs_1[31]~q ;
wire \io_w_dmem_dat_data[31]~47_combout ;

wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a31_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a31_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a0_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a4_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a3_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a2_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a1_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a24_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a23_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a23_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a24_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a22_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a22_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a21_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a21_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a20_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a19_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a19_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a20_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a18_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a18_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a17_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a17_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a16_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a15_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a16_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a14_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a13_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a28_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a28_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a30_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a30_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a29_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a27_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a27_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a29_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a26_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a26_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a25_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a25_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a12_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a11_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a10_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a9_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a8_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a7_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a6_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus ;
wire [143:0] \_T_3543_rtl_1|auto_generated|ram_block1a5_PORTBDATAOUT_bus ;

assign \_T_3543_rtl_1|auto_generated|ram_block1a31~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a31_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a31~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a31_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a0~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a0~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a0_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a4~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a4_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a3~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a3_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a3~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a4~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a2~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a2_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a2~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a1~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a1_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a1~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a24~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a24_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a23~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a23_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a23~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a23_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a24~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a24_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a22~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a22_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a22~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a22_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a21~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a21_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a21~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a21_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a20~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a20_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a19~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a19_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a19~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a19_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a20~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a20_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a18~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a18_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a18~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a18_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a17~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a17_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a17~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a17_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a16~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a16_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a15~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a15_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a15~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a16~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a16_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a14~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a14_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a14~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a13~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a13~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a13_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a28~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a28_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a28~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a28_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a30~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a30_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a30~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a30_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a29~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a29_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a27~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a27_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a27~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a27_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a29~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a29_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a26~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a26_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a26~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a26_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a25~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a25_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a25~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a25_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a12~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a12_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a11~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a11_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a11~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a12~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a10~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a10_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a10~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a9~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a9~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a9_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a8~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a8_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a7~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a7_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a7~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a8~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a6~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a6_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a6~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_0|auto_generated|ram_block1a5~portbdataout  = \_T_3543_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus [0];

assign \_T_3543_rtl_1|auto_generated|ram_block1a5~portbdataout  = \_T_3543_rtl_1|auto_generated|ram_block1a5_PORTBDATAOUT_bus [0];

kyogenrv_fpga_ALU alu(
	.ex_ctrl_alu_op1_0(\ex_ctrl_alu_op1[0]~q ),
	.ex_ctrl_alu_op1_1(\ex_ctrl_alu_op1[1]~q ),
	.ex_ctrl_imm_type011(\ex_ctrl_imm_type.011~q ),
	.ex_ctrl_alu_func_0(\ex_ctrl_alu_func[0]~q ),
	._T_3_0(\alu|_T_3[0]~0_combout ),
	._T_3_1(\alu|_T_3[1]~2_combout ),
	._T_3_2(\alu|_T_3[2]~4_combout ),
	._T_3_3(\alu|_T_3[3]~6_combout ),
	._T_3_4(\alu|_T_3[4]~8_combout ),
	._T_3_5(\alu|_T_3[5]~10_combout ),
	._T_3_6(\alu|_T_3[6]~12_combout ),
	._T_3_7(\alu|_T_3[7]~14_combout ),
	._T_3_8(\alu|_T_3[8]~16_combout ),
	._T_3_9(\alu|_T_3[9]~18_combout ),
	._T_3_10(\alu|_T_3[10]~20_combout ),
	._T_3_11(\alu|_T_3[11]~22_combout ),
	._T_3_12(\alu|_T_3[12]~24_combout ),
	._T_3_13(\alu|_T_3[13]~26_combout ),
	._T_3_14(\alu|_T_3[14]~28_combout ),
	._T_3_15(\alu|_T_3[15]~30_combout ),
	._T_3_16(\alu|_T_3[16]~32_combout ),
	._T_3_17(\alu|_T_3[17]~34_combout ),
	._T_3_18(\alu|_T_3[18]~36_combout ),
	._T_3_19(\alu|_T_3[19]~38_combout ),
	._T_3_20(\alu|_T_3[20]~40_combout ),
	._T_3_21(\alu|_T_3[21]~42_combout ),
	._T_3_22(\alu|_T_3[22]~44_combout ),
	._T_3_23(\alu|_T_3[23]~46_combout ),
	._T_3_24(\alu|_T_3[24]~48_combout ),
	._T_3_25(\alu|_T_3[25]~50_combout ),
	._T_3_26(\alu|_T_3[26]~52_combout ),
	._T_3_27(\alu|_T_3[27]~54_combout ),
	._T_3_28(\alu|_T_3[28]~56_combout ),
	._T_3_29(\alu|_T_3[29]~58_combout ),
	._T_3_30(\alu|_T_3[30]~60_combout ),
	._T_3_31(\alu|_T_3[31]~62_combout ),
	.csr_io_alu_op1_0(\csr_io_alu_op1[0]~4_combout ),
	.ex_ctrl_alu_op201(\ex_ctrl_alu_op2.01~q ),
	.ex_ctrl_alu_op210(\ex_ctrl_alu_op2.10~q ),
	.csr_io_alu_op2_1(\csr_io_alu_op2[1]~0_combout ),
	.ex_reg_rs2_bypass_1(\ex_reg_rs2_bypass[1]~9_combout ),
	.io_sw_r_ex_imm_1(\io_sw_r_ex_imm[1]~1_combout ),
	.csr_io_alu_op2_11(\csr_io_alu_op2[1]~1_combout ),
	.csr_io_alu_op2_0(\csr_io_alu_op2[0]~2_combout ),
	.alu_io_op2_3(\alu_io_op2[3]~42_combout ),
	.ex_reg_rs2_bypass_0(\ex_reg_rs2_bypass[0]~11_combout ),
	._T_3681(\_T_3681~3_combout ),
	.ex_reg_rs2_bypass_01(\ex_reg_rs2_bypass[0]~14_combout ),
	.csr_io_alu_op2_01(\csr_io_alu_op2[0]~3_combout ),
	._T_123_31(\alu|_T_123[31]~combout ),
	.alu_io_op2_9(\alu_io_op2[9]~45_combout ),
	.alu_io_op2_8(\alu_io_op2[8]~47_combout ),
	.alu_io_op2_10(\alu_io_op2[10]~49_combout ),
	.alu_io_op2_11(\alu_io_op2[11]~51_combout ),
	._T_123_11(\alu|_T_123[11]~combout ),
	.mem_csr_data_12(\mem_csr_data[12]~q ),
	.mem_csr_data_13(\mem_csr_data[13]~q ),
	.alu_io_op2_13(\alu_io_op2[13]~52_combout ),
	.ex_reg_rs2_bypass_13(\ex_reg_rs2_bypass[13]~45_combout ),
	.ex_reg_rs2_bypass_131(\ex_reg_rs2_bypass[13]~46_combout ),
	.alu_io_op2_12(\alu_io_op2[12]~53_combout ),
	.ex_reg_rs2_bypass_12(\ex_reg_rs2_bypass[12]~49_combout ),
	.mem_csr_data_14(\mem_csr_data[14]~q ),
	.alu_io_op2_14(\alu_io_op2[14]~54_combout ),
	.ex_reg_rs2_bypass_14(\ex_reg_rs2_bypass[14]~53_combout ),
	.ex_reg_rs2_bypass_15(\ex_reg_rs2_bypass[15]~58_combout ),
	.alu_io_op2_15(\alu_io_op2[15]~55_combout ),
	._T_123_15(\alu|_T_123[15]~combout ),
	.alu_io_op2_17(\alu_io_op2[17]~56_combout ),
	.ex_reg_rs2_bypass_17(\ex_reg_rs2_bypass[17]~62_combout ),
	.alu_io_op2_16(\alu_io_op2[16]~57_combout ),
	.ex_reg_rs2_bypass_16(\ex_reg_rs2_bypass[16]~66_combout ),
	.alu_io_op2_18(\alu_io_op2[18]~58_combout ),
	.ex_reg_rs2_bypass_18(\ex_reg_rs2_bypass[18]~70_combout ),
	.ex_reg_rs2_bypass_19(\ex_reg_rs2_bypass[19]~74_combout ),
	.alu_io_op2_19(\alu_io_op2[19]~59_combout ),
	._T_123_19(\alu|_T_123[19]~combout ),
	.alu_io_op2_4(\alu_io_op2[4]~61_combout ),
	.io_sw_r_ex_imm_4(\io_sw_r_ex_imm[4]~4_combout ),
	.alu_io_op2_41(\alu_io_op2[4]~62_combout ),
	.ex_ctrl_alu_func_3(\ex_ctrl_alu_func[3]~q ),
	.alu_io_op2_2(\alu_io_op2[2]~63_combout ),
	._T_123_2(\alu|_T_123[2]~combout ),
	.alu_io_op2_31(\alu_io_op2[3]~65_combout ),
	.io_sw_r_ex_imm_3(\io_sw_r_ex_imm[3]~8_combout ),
	.alu_io_op2_32(\alu_io_op2[3]~66_combout ),
	.alu_io_op2_5(\alu_io_op2[5]~68_combout ),
	.alu_io_op2_6(\alu_io_op2[6]~70_combout ),
	.alu_io_op2_7(\alu_io_op2[7]~72_combout ),
	._T_123_7(\alu|_T_123[7]~combout ),
	.alu_io_op1_23(\alu_io_op1[23]~60_combout ),
	.alu_io_op1_27(\alu_io_op1[27]~61_combout ),
	.ex_ctrl_alu_func_1(\ex_ctrl_alu_func[1]~q ),
	.ex_ctrl_alu_func_2(\ex_ctrl_alu_func[2]~q ),
	.LessThan0(\alu|LessThan0~0_combout ),
	._T_125(\alu|_T_125~20_combout ),
	.alu_io_op1_31(\alu_io_op1[31]~62_combout ),
	.csr_io_alu_op1_01(\csr_io_alu_op1[0]~5_combout ),
	.alu_io_op1_30(\alu_io_op1[30]~63_combout ),
	.csr_io_alu_op1_1(\csr_io_alu_op1[1]~6_combout ),
	.ShiftRight0(\alu|ShiftRight0~38_combout ),
	.alu_io_op1_8(\alu_io_op1[8]~64_combout ),
	.alu_io_op1_7(\alu_io_op1[7]~65_combout ),
	.alu_io_op1_24(\alu_io_op1[24]~66_combout ),
	.alu_io_op1_4(\alu_io_op1[4]~67_combout ),
	.alu_io_op1_3(\alu_io_op1[3]~68_combout ),
	.alu_io_op1_28(\alu_io_op1[28]~69_combout ),
	.alu_io_op1_6(\alu_io_op1[6]~70_combout ),
	.alu_io_op1_25(\alu_io_op1[25]~71_combout ),
	.alu_io_op1_5(\alu_io_op1[5]~72_combout ),
	.alu_io_op1_26(\alu_io_op1[26]~73_combout ),
	.alu_io_op1_2(\alu_io_op1[2]~74_combout ),
	.alu_io_op1_29(\alu_io_op1[29]~75_combout ),
	.alu_io_op1_12(\alu_io_op1[12]~76_combout ),
	.alu_io_op1_19(\alu_io_op1[19]~77_combout ),
	.alu_io_op1_11(\alu_io_op1[11]~78_combout ),
	.alu_io_op1_20(\alu_io_op1[20]~79_combout ),
	.alu_io_op1_10(\alu_io_op1[10]~80_combout ),
	.alu_io_op1_21(\alu_io_op1[21]~81_combout ),
	.alu_io_op1_9(\alu_io_op1[9]~82_combout ),
	.alu_io_op1_22(\alu_io_op1[22]~83_combout ),
	.alu_io_op1_16(\alu_io_op1[16]~84_combout ),
	.alu_io_op1_15(\alu_io_op1[15]~85_combout ),
	.alu_io_op1_14(\alu_io_op1[14]~86_combout ),
	.alu_io_op1_17(\alu_io_op1[17]~87_combout ),
	.alu_io_op1_13(\alu_io_op1[13]~88_combout ),
	.alu_io_op1_18(\alu_io_op1[18]~89_combout ),
	.ShiftRight01(\alu|ShiftRight0~94_combout ),
	.ShiftRight02(\alu|ShiftRight0~126_combout ),
	.ShiftRight03(\alu|ShiftRight0~128_combout ),
	.io_out_0(\alu|io_out[0]~1_combout ),
	.ShiftRight04(\alu|ShiftRight0~130_combout ),
	.ShiftRight05(\alu|ShiftRight0~150_combout ),
	.ShiftRight06(\alu|ShiftRight0~152_combout ),
	.ShiftRight07(\alu|ShiftRight0~167_combout ),
	.ShiftRight08(\alu|ShiftRight0~173_combout ),
	.ShiftRight09(\alu|ShiftRight0~175_combout ),
	.ShiftRight010(\alu|ShiftRight0~180_combout ),
	.ShiftRight011(\alu|ShiftRight0~183_combout ),
	.ShiftRight012(\alu|ShiftRight0~188_combout ),
	.ShiftRight013(\alu|ShiftRight0~190_combout ),
	.ShiftRight014(\alu|ShiftRight0~195_combout ),
	.ShiftRight015(\alu|ShiftRight0~197_combout ),
	.ShiftRight016(\alu|ShiftRight0~198_combout ),
	.ShiftRight017(\alu|ShiftRight0~203_combout ),
	._T_123_13(\alu|_T_123[13]~combout ),
	.ShiftRight018(\alu|ShiftRight0~209_combout ),
	.ShiftRight019(\alu|ShiftRight0~216_combout ),
	.ShiftRight020(\alu|ShiftRight0~217_combout ),
	.ShiftRight021(\alu|ShiftRight0~222_combout ),
	._T_139_18(\alu|_T_139[18]~combout ),
	.ShiftRight022(\alu|ShiftRight0~228_combout ),
	.ShiftRight023(\alu|ShiftRight0~233_combout ),
	.ShiftRight024(\alu|ShiftRight0~236_combout ),
	.ShiftRight025(\alu|ShiftRight0~240_combout ),
	.csr_io_alu_op1_11(\csr_io_alu_op1[1]~7_combout ),
	.csr_io_alu_op1_02(\csr_io_alu_op1[0]~8_combout ),
	.alu_io_op1_281(\alu_io_op1[28]~90_combout ),
	.alu_io_op1_291(\alu_io_op1[29]~91_combout ),
	.alu_io_op2_29(\alu_io_op2[29]~73_combout ),
	.alu_io_op2_28(\alu_io_op2[28]~74_combout ),
	.alu_io_op1_301(\alu_io_op1[30]~92_combout ),
	.alu_io_op2_30(\alu_io_op2[30]~75_combout ),
	.alu_io_op1_311(\alu_io_op1[31]~93_combout ),
	.alu_io_op2_311(\alu_io_op2[31]~76_combout ),
	.alu_io_op1_81(\alu_io_op1[8]~94_combout ),
	.alu_io_op1_91(\alu_io_op1[9]~95_combout ),
	.alu_io_op1_101(\alu_io_op1[10]~96_combout ),
	.alu_io_op1_111(\alu_io_op1[11]~97_combout ),
	.alu_io_op1_121(\alu_io_op1[12]~98_combout ),
	.alu_io_op1_131(\alu_io_op1[13]~99_combout ),
	.alu_io_op2_131(\alu_io_op2[13]~77_combout ),
	.alu_io_op2_121(\alu_io_op2[12]~78_combout ),
	.alu_io_op1_141(\alu_io_op1[14]~100_combout ),
	.alu_io_op2_141(\alu_io_op2[14]~79_combout ),
	.alu_io_op1_151(\alu_io_op1[15]~101_combout ),
	.alu_io_op1_161(\alu_io_op1[16]~102_combout ),
	.alu_io_op1_171(\alu_io_op1[17]~103_combout ),
	.alu_io_op2_171(\alu_io_op2[17]~80_combout ),
	.alu_io_op2_161(\alu_io_op2[16]~81_combout ),
	.alu_io_op1_181(\alu_io_op1[18]~104_combout ),
	.alu_io_op2_181(\alu_io_op2[18]~82_combout ),
	.alu_io_op1_191(\alu_io_op1[19]~105_combout ),
	.alu_io_op1_41(\alu_io_op1[4]~106_combout ),
	.alu_io_op1_210(\alu_io_op1[2]~107_combout ),
	.alu_io_op1_51(\alu_io_op1[5]~108_combout ),
	.alu_io_op1_32(\alu_io_op1[3]~109_combout ),
	.alu_io_op1_61(\alu_io_op1[6]~110_combout ),
	.alu_io_op1_71(\alu_io_op1[7]~111_combout ),
	.alu_io_op1_201(\alu_io_op1[20]~112_combout ),
	.alu_io_op1_211(\alu_io_op1[21]~113_combout ),
	.alu_io_op2_21(\alu_io_op2[21]~83_combout ),
	.alu_io_op2_20(\alu_io_op2[20]~84_combout ),
	.alu_io_op1_221(\alu_io_op1[22]~114_combout ),
	.alu_io_op2_22(\alu_io_op2[22]~85_combout ),
	.alu_io_op2_23(\alu_io_op2[23]~86_combout ),
	._T_123_23(\alu|_T_123[23]~combout ),
	.alu_io_op1_241(\alu_io_op1[24]~115_combout ),
	.alu_io_op1_251(\alu_io_op1[25]~116_combout ),
	.alu_io_op2_25(\alu_io_op2[25]~87_combout ),
	.alu_io_op2_24(\alu_io_op2[24]~88_combout ),
	.alu_io_op1_261(\alu_io_op1[26]~117_combout ),
	.alu_io_op2_26(\alu_io_op2[26]~89_combout ),
	.alu_io_op2_27(\alu_io_op2[27]~90_combout ),
	._T_123_27(\alu|_T_123[27]~combout ),
	.alu_io_op1_271(\alu_io_op1[27]~118_combout ),
	.alu_io_op1_231(\alu_io_op1[23]~119_combout ),
	.alu_io_op2_210(\alu_io_op2[2]~91_combout ),
	._T_123_29(\alu|_T_123[29]~combout ),
	.ShiftRight026(\alu|ShiftRight0~249_combout ),
	.ShiftRight027(\alu|ShiftRight0~250_combout ),
	._T_123_17(\alu|_T_123[17]~combout ),
	.ShiftRight028(\alu|ShiftRight0~251_combout ),
	.ShiftRight029(\alu|ShiftRight0~253_combout ),
	.ShiftRight030(\alu|ShiftRight0~254_combout ),
	.ShiftRight031(\alu|ShiftRight0~256_combout ),
	._T_123_21(\alu|_T_123[21]~combout ),
	._T_123_25(\alu|_T_123[25]~combout ));

kyogenrv_fpga_CSR csr(
	.ex_j_check(\ex_j_check~q ),
	.ex_ctrl_mem_wr01(\ex_ctrl_mem_wr.01~q ),
	._T_3549(\_T_3549~q ),
	.mepc_2(\csr|mepc[2]~q ),
	.mepc_3(\csr|mepc[3]~q ),
	.mepc_4(\csr|mepc[4]~q ),
	.mepc_5(\csr|mepc[5]~q ),
	.mepc_6(\csr|mepc[6]~q ),
	.mepc_7(\csr|mepc[7]~q ),
	.mepc_8(\csr|mepc[8]~q ),
	.mepc_9(\csr|mepc[9]~q ),
	.mepc_10(\csr|mepc[10]~q ),
	.mepc_11(\csr|mepc[11]~q ),
	.mepc_12(\csr|mepc[12]~q ),
	.mepc_13(\csr|mepc[13]~q ),
	.mepc_14(\csr|mepc[14]~q ),
	.mepc_15(\csr|mepc[15]~q ),
	.mepc_16(\csr|mepc[16]~q ),
	.mepc_17(\csr|mepc[17]~q ),
	.mepc_18(\csr|mepc[18]~q ),
	.mepc_19(\csr|mepc[19]~q ),
	.mepc_20(\csr|mepc[20]~q ),
	.mepc_21(\csr|mepc[21]~q ),
	.mepc_22(\csr|mepc[22]~q ),
	.mepc_23(\csr|mepc[23]~q ),
	.mepc_24(\csr|mepc[24]~q ),
	.mepc_25(\csr|mepc[25]~q ),
	.mepc_26(\csr|mepc[26]~q ),
	.mepc_27(\csr|mepc[27]~q ),
	.mepc_28(\csr|mepc[28]~q ),
	.mepc_29(\csr|mepc[29]~q ),
	.mepc_30(\csr|mepc[30]~q ),
	.mepc_31(\csr|mepc[31]~q ),
	.ex_b_check(\ex_b_check~q ),
	.inst_kill(\inst_kill~0_combout ),
	.ex_npc_0(\ex_npc[0]~q ),
	.ex_npc_1(\ex_npc[1]~q ),
	.Equal56(\Equal56~0_combout ),
	.ex_pc_4(\ex_pc[4]~q ),
	.ex_pc_5(\ex_pc[5]~q ),
	.ex_pc_6(\ex_pc[6]~q ),
	.ex_pc_7(\ex_pc[7]~q ),
	.ex_pc_2(\ex_pc[2]~q ),
	.ex_pc_3(\ex_pc[3]~q ),
	.ex_pc_8(\ex_pc[8]~q ),
	.ex_pc_9(\ex_pc[9]~q ),
	.ex_pc_10(\ex_pc[10]~q ),
	.ex_pc_11(\ex_pc[11]~q ),
	.ex_pc_12(\ex_pc[12]~q ),
	.ex_pc_13(\ex_pc[13]~q ),
	.ex_pc_14(\ex_pc[14]~q ),
	.ex_pc_15(\ex_pc[15]~q ),
	.ex_pc_16(\ex_pc[16]~q ),
	.ex_pc_17(\ex_pc[17]~q ),
	.ex_pc_18(\ex_pc[18]~q ),
	.ex_pc_19(\ex_pc[19]~q ),
	.ex_pc_20(\ex_pc[20]~q ),
	.ex_pc_21(\ex_pc[21]~q ),
	.ex_pc_22(\ex_pc[22]~q ),
	.ex_pc_23(\ex_pc[23]~q ),
	.ex_pc_24(\ex_pc[24]~q ),
	.ex_pc_25(\ex_pc[25]~q ),
	.ex_pc_26(\ex_pc[26]~q ),
	.ex_pc_27(\ex_pc[27]~q ),
	.ex_pc_28(\ex_pc[28]~q ),
	.ex_pc_29(\ex_pc[29]~q ),
	.ex_pc_30(\ex_pc[30]~q ),
	.ex_pc_31(\ex_pc[31]~q ),
	.Equal561(\Equal56~10_combout ),
	.ex_ctrl_legal(\ex_ctrl_legal~q ),
	.Equal59(\Equal59~1_combout ),
	.ex_csr_addr_0(\ex_csr_addr[0]~q ),
	.ex_csr_addr_1(\ex_csr_addr[1]~q ),
	.ex_csr_addr_2(\ex_csr_addr[2]~q ),
	.ex_csr_addr_3(\ex_csr_addr[3]~q ),
	.ex_csr_addr_4(\ex_csr_addr[4]~q ),
	.Equal62(\Equal62~0_combout ),
	.ex_inst_8(\ex_inst[8]~q ),
	.ex_ctrl_imm_type001(\ex_ctrl_imm_type.001~q ),
	.csr_io_alu_op2_1(\csr_io_alu_op2[1]~1_combout ),
	.ex_inst_7(\ex_inst[7]~q ),
	.csr_io_alu_op2_0(\csr_io_alu_op2[0]~3_combout ),
	.ex_ctrl_mask_type_0(\ex_ctrl_mask_type[0]~q ),
	.ex_ctrl_mask_type_2(\ex_ctrl_mask_type[2]~q ),
	.ex_ctrl_mask_type_1(\ex_ctrl_mask_type[1]~q ),
	.io_expt1(\csr|io_expt~0_combout ),
	.waitrequest_reset_override(waitrequest_reset_override),
	.wait_latency_counter_0(wait_latency_counter_0),
	.mem_ctrl_mem_wr10(mem_ctrl_mem_wr10),
	.wait_latency_counter_1(wait_latency_counter_1),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.ex_inst_9(\ex_inst[9]~q ),
	.ex_inst_10(\ex_inst[10]~q ),
	.ex_inst_11(\ex_inst[11]~q ),
	._T_3557(\_T_3557~6_combout ),
	.mcause_0(\csr|mcause[0]~6_combout ),
	.ex_csr_cmd_2(\ex_csr_cmd[2]~q ),
	.ex_csr_cmd_0(\ex_csr_cmd[0]~q ),
	.ex_csr_cmd_1(\ex_csr_cmd[1]~q ),
	.ex_csr_addr_8(\ex_csr_addr[8]~q ),
	.isEcall(\csr|isEcall~0_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.mepc_0(\csr|mepc[0]~q ),
	.io_expt2(\csr|io_expt~combout ),
	.mtvec_0(\csr|mtvec[0]~q ),
	.ex_csr_addr_9(\ex_csr_addr[9]~q ),
	.ex_csr_addr_11(\ex_csr_addr[11]~q ),
	.ex_csr_addr_10(\ex_csr_addr[10]~q ),
	.ex_inst_13(\ex_inst[13]~q ),
	.ex_inst_12(\ex_inst[12]~q ),
	.ex_inst_14(\ex_inst[14]~q ),
	.ex_csr_addr_5(\ex_csr_addr[5]~q ),
	.ex_csr_addr_6(\ex_csr_addr[6]~q ),
	.ex_csr_addr_7(\ex_csr_addr[7]~q ),
	.mepc_1(\csr|mepc[1]~q ),
	.mtvec_1(\csr|mtvec[1]~q ),
	.io_out_1(\csr|io_out[1]~16_combout ),
	.io_out_0(\csr|io_out[0]~24_combout ),
	.mtvec_2(\csr|mtvec[2]~q ),
	.mtvec_3(\csr|mtvec[3]~q ),
	.mtvec_4(\csr|mtvec[4]~q ),
	.mtvec_5(\csr|mtvec[5]~q ),
	.mtvec_6(\csr|mtvec[6]~q ),
	.mtvec_7(\csr|mtvec[7]~q ),
	.mtvec_8(\csr|mtvec[8]~q ),
	.mtvec_9(\csr|mtvec[9]~q ),
	.mtvec_10(\csr|mtvec[10]~q ),
	.mtvec_11(\csr|mtvec[11]~q ),
	.mtvec_12(\csr|mtvec[12]~q ),
	.mtvec_13(\csr|mtvec[13]~q ),
	.mtvec_14(\csr|mtvec[14]~q ),
	.mtvec_15(\csr|mtvec[15]~q ),
	.mtvec_16(\csr|mtvec[16]~q ),
	.mtvec_17(\csr|mtvec[17]~q ),
	.mtvec_18(\csr|mtvec[18]~q ),
	.mtvec_19(\csr|mtvec[19]~q ),
	.mtvec_20(\csr|mtvec[20]~q ),
	.mtvec_21(\csr|mtvec[21]~q ),
	.mtvec_22(\csr|mtvec[22]~q ),
	.mtvec_23(\csr|mtvec[23]~q ),
	.mtvec_24(\csr|mtvec[24]~q ),
	.mtvec_25(\csr|mtvec[25]~q ),
	.mtvec_26(\csr|mtvec[26]~q ),
	.mtvec_27(\csr|mtvec[27]~q ),
	.mtvec_28(\csr|mtvec[28]~q ),
	.mtvec_29(\csr|mtvec[29]~q ),
	.mtvec_30(\csr|mtvec[30]~q ),
	.mtvec_31(\csr|mtvec[31]~q ),
	.csr_io_in_0(\csr_io_in[0]~6_combout ),
	.io_out_28(\csr|io_out[28]~31_combout ),
	.io_out_29(\csr|io_out[29]~36_combout ),
	.io_out_291(\csr|io_out[29]~37_combout ),
	.io_out_30(\csr|io_out[30]~45_combout ),
	.io_out_31(\csr|io_out[31]~52_combout ),
	.io_out_8(\csr|io_out[8]~59_combout ),
	.io_out_9(\csr|io_out[9]~66_combout ),
	.io_out_10(\csr|io_out[10]~72_combout ),
	.io_out_11(\csr|io_out[11]~79_combout ),
	.io_out_12(\csr|io_out[12]~86_combout ),
	.io_out_13(\csr|io_out[13]~93_combout ),
	.io_out_14(\csr|io_out[14]~100_combout ),
	.io_out_15(\csr|io_out[15]~107_combout ),
	.io_out_16(\csr|io_out[16]~114_combout ),
	.io_out_17(\csr|io_out[17]~121_combout ),
	.io_out_18(\csr|io_out[18]~128_combout ),
	.io_out_19(\csr|io_out[19]~135_combout ),
	.io_out_4(\csr|io_out[4]~142_combout ),
	.io_out_2(\csr|io_out[2]~150_combout ),
	.io_out_3(\csr|io_out[3]~159_combout ),
	.io_out_5(\csr|io_out[5]~166_combout ),
	.io_out_6(\csr|io_out[6]~173_combout ),
	.io_out_7(\csr|io_out[7]~181_combout ),
	.io_out_20(\csr|io_out[20]~188_combout ),
	.io_out_21(\csr|io_out[21]~193_combout ),
	.io_out_211(\csr|io_out[21]~194_combout ),
	.io_out_22(\csr|io_out[22]~202_combout ),
	.io_out_23(\csr|io_out[23]~209_combout ),
	.io_out_24(\csr|io_out[24]~216_combout ),
	.io_out_25(\csr|io_out[25]~221_combout ),
	.io_out_251(\csr|io_out[25]~222_combout ),
	.io_out_26(\csr|io_out[26]~230_combout ),
	.io_out_27(\csr|io_out[27]~235_combout ),
	.io_out_271(\csr|io_out[27]~236_combout ),
	.csr_io_in_1(\csr_io_in[1]~10_combout ),
	.ex_inst_0(\ex_inst[0]~q ),
	.ex_inst_1(\ex_inst[1]~q ),
	.ex_inst_4(\ex_inst[4]~q ),
	.ex_inst_2(\ex_inst[2]~q ),
	.ex_inst_3(\ex_inst[3]~q ),
	.ex_inst_5(\ex_inst[5]~q ),
	.ex_inst_6(\ex_inst[6]~q ),
	.csr_io_in_2(\csr_io_in[2]~14_combout ),
	.csr_io_in_3(\csr_io_in[3]~18_combout ),
	.csr_io_in_4(\csr_io_in[4]~22_combout ),
	.csr_io_in_5(\csr_io_in[5]~25_combout ),
	.csr_io_in_6(\csr_io_in[6]~28_combout ),
	.csr_io_in_7(\csr_io_in[7]~31_combout ),
	.csr_io_in_8(\csr_io_in[8]~34_combout ),
	.csr_io_in_9(\csr_io_in[9]~37_combout ),
	.csr_io_in_10(\csr_io_in[10]~40_combout ),
	.csr_io_in_11(\csr_io_in[11]~43_combout ),
	.csr_io_in_12(\csr_io_in[12]~46_combout ),
	.csr_io_in_13(\csr_io_in[13]~49_combout ),
	.csr_io_in_14(\csr_io_in[14]~52_combout ),
	.csr_io_in_15(\csr_io_in[15]~55_combout ),
	.csr_io_in_16(\csr_io_in[16]~58_combout ),
	.csr_io_in_17(\csr_io_in[17]~61_combout ),
	.csr_io_in_18(\csr_io_in[18]~64_combout ),
	.csr_io_in_19(\csr_io_in[19]~67_combout ),
	.csr_io_in_20(\csr_io_in[20]~70_combout ),
	.csr_io_in_21(\csr_io_in[21]~73_combout ),
	.csr_io_in_22(\csr_io_in[22]~76_combout ),
	.csr_io_in_23(\csr_io_in[23]~79_combout ),
	.csr_io_in_24(\csr_io_in[24]~82_combout ),
	.csr_io_in_25(\csr_io_in[25]~85_combout ),
	.csr_io_in_26(\csr_io_in[26]~88_combout ),
	.csr_io_in_27(\csr_io_in[27]~91_combout ),
	.csr_io_in_28(\csr_io_in[28]~94_combout ),
	.csr_io_in_29(\csr_io_in[29]~97_combout ),
	.csr_io_in_30(\csr_io_in[30]~100_combout ),
	.csr_io_in_31(\csr_io_in[31]~104_combout ),
	.csr_io_alu_op1_1(\csr_io_alu_op1[1]~7_combout ),
	.csr_io_alu_op1_0(\csr_io_alu_op1[0]~8_combout ),
	.clock(clk_clk));

dffeas ex_j_check(
	.clk(clk_clk),
	.d(\_GEN_32~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_j_check~q ),
	.prn(vcc));
defparam ex_j_check.is_wysiwyg = "true";
defparam ex_j_check.power_up = "low";

dffeas _T_3549(
	.clk(!clk_clk),
	.d(\_GEN_9~combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(\_T_3549~q ),
	.prn(vcc));
defparam _T_3549.is_wysiwyg = "true";
defparam _T_3549.power_up = "low";

dffeas ex_b_check(
	.clk(clk_clk),
	.d(\_GEN_33~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_b_check~q ),
	.prn(vcc));
defparam ex_b_check.is_wysiwyg = "true";
defparam ex_b_check.power_up = "low";

cyclone10lp_lcell_comb \Equal56~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\ex_npc[0]~q ),
	.datad(\ex_npc[1]~q ),
	.cin(gnd),
	.combout(\Equal56~0_combout ),
	.cout());
defparam \Equal56~0 .lut_mask = 16'h000F;
defparam \Equal56~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal56~1 (
	.dataa(\ex_pc[4]~q ),
	.datab(\ex_pc[5]~q ),
	.datac(\ex_pc[6]~q ),
	.datad(\ex_pc[7]~q ),
	.cin(gnd),
	.combout(\Equal56~1_combout ),
	.cout());
defparam \Equal56~1 .lut_mask = 16'h0001;
defparam \Equal56~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal56~2 (
	.dataa(\Equal56~0_combout ),
	.datab(\Equal56~1_combout ),
	.datac(\ex_pc[2]~q ),
	.datad(\ex_pc[3]~q ),
	.cin(gnd),
	.combout(\Equal56~2_combout ),
	.cout());
defparam \Equal56~2 .lut_mask = 16'h0008;
defparam \Equal56~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal56~3 (
	.dataa(\ex_pc[8]~q ),
	.datab(\ex_pc[9]~q ),
	.datac(\ex_pc[10]~q ),
	.datad(\ex_pc[11]~q ),
	.cin(gnd),
	.combout(\Equal56~3_combout ),
	.cout());
defparam \Equal56~3 .lut_mask = 16'h0001;
defparam \Equal56~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal56~4 (
	.dataa(\ex_pc[12]~q ),
	.datab(\ex_pc[13]~q ),
	.datac(\ex_pc[14]~q ),
	.datad(\ex_pc[15]~q ),
	.cin(gnd),
	.combout(\Equal56~4_combout ),
	.cout());
defparam \Equal56~4 .lut_mask = 16'h0001;
defparam \Equal56~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal56~5 (
	.dataa(\ex_pc[16]~q ),
	.datab(\ex_pc[17]~q ),
	.datac(\ex_pc[18]~q ),
	.datad(\ex_pc[19]~q ),
	.cin(gnd),
	.combout(\Equal56~5_combout ),
	.cout());
defparam \Equal56~5 .lut_mask = 16'h0001;
defparam \Equal56~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal56~6 (
	.dataa(\ex_pc[20]~q ),
	.datab(\ex_pc[21]~q ),
	.datac(\ex_pc[22]~q ),
	.datad(\ex_pc[23]~q ),
	.cin(gnd),
	.combout(\Equal56~6_combout ),
	.cout());
defparam \Equal56~6 .lut_mask = 16'h0001;
defparam \Equal56~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal56~7 (
	.dataa(\ex_pc[24]~q ),
	.datab(\ex_pc[25]~q ),
	.datac(\ex_pc[26]~q ),
	.datad(\ex_pc[27]~q ),
	.cin(gnd),
	.combout(\Equal56~7_combout ),
	.cout());
defparam \Equal56~7 .lut_mask = 16'h0001;
defparam \Equal56~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal56~8 (
	.dataa(\ex_pc[28]~q ),
	.datab(\ex_pc[29]~q ),
	.datac(\ex_pc[30]~q ),
	.datad(\ex_pc[31]~q ),
	.cin(gnd),
	.combout(\Equal56~8_combout ),
	.cout());
defparam \Equal56~8 .lut_mask = 16'h0001;
defparam \Equal56~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal56~9 (
	.dataa(\Equal56~5_combout ),
	.datab(\Equal56~6_combout ),
	.datac(\Equal56~7_combout ),
	.datad(\Equal56~8_combout ),
	.cin(gnd),
	.combout(\Equal56~9_combout ),
	.cout());
defparam \Equal56~9 .lut_mask = 16'h8000;
defparam \Equal56~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal56~10 (
	.dataa(\Equal56~2_combout ),
	.datab(\Equal56~3_combout ),
	.datac(\Equal56~4_combout ),
	.datad(\Equal56~9_combout ),
	.cin(gnd),
	.combout(\Equal56~10_combout ),
	.cout());
defparam \Equal56~10 .lut_mask = 16'h8000;
defparam \Equal56~10 .sum_lutc_input = "datac";

dffeas ex_ctrl_legal(
	.clk(clk_clk),
	.d(\ex_ctrl_legal~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_legal~q ),
	.prn(vcc));
defparam ex_ctrl_legal.is_wysiwyg = "true";
defparam ex_ctrl_legal.power_up = "low";

cyclone10lp_lcell_comb \csr_io_alu_op1[0]~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\ex_ctrl_alu_op1[0]~q ),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\csr_io_alu_op1[0]~4_combout ),
	.cout());
defparam \csr_io_alu_op1[0]~4 .lut_mask = 16'h0FF0;
defparam \csr_io_alu_op1[0]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3557~0 (
	.dataa(\ex_inst[7]~q ),
	.datab(\ex_inst[8]~q ),
	.datac(\id_inst[16]~q ),
	.datad(\id_inst[15]~q ),
	.cin(gnd),
	.combout(\_T_3557~0_combout ),
	.cout());
defparam \_T_3557~0 .lut_mask = 16'h8241;
defparam \_T_3557~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3557~1 (
	.dataa(\ex_inst[9]~q ),
	.datab(\ex_inst[10]~q ),
	.datac(\id_inst[18]~q ),
	.datad(\id_inst[17]~q ),
	.cin(gnd),
	.combout(\_T_3557~1_combout ),
	.cout());
defparam \_T_3557~1 .lut_mask = 16'h8241;
defparam \_T_3557~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3557~2 (
	.dataa(\_T_3557~0_combout ),
	.datab(\_T_3557~1_combout ),
	.datac(\ex_inst[11]~q ),
	.datad(\id_inst[19]~q ),
	.cin(gnd),
	.combout(\_T_3557~2_combout ),
	.cout());
defparam \_T_3557~2 .lut_mask = 16'h8008;
defparam \_T_3557~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3557~3 (
	.dataa(\ex_inst[7]~q ),
	.datab(\ex_inst[8]~q ),
	.datac(\id_inst[21]~q ),
	.datad(\id_inst[20]~q ),
	.cin(gnd),
	.combout(\_T_3557~3_combout ),
	.cout());
defparam \_T_3557~3 .lut_mask = 16'h8241;
defparam \_T_3557~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3557~4 (
	.dataa(\ex_inst[9]~q ),
	.datab(\ex_inst[10]~q ),
	.datac(\id_inst[23]~q ),
	.datad(\id_inst[22]~q ),
	.cin(gnd),
	.combout(\_T_3557~4_combout ),
	.cout());
defparam \_T_3557~4 .lut_mask = 16'h8241;
defparam \_T_3557~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3557~5 (
	.dataa(\_T_3557~3_combout ),
	.datab(\_T_3557~4_combout ),
	.datac(\ex_inst[11]~q ),
	.datad(\id_inst[24]~q ),
	.cin(gnd),
	.combout(\_T_3557~5_combout ),
	.cout());
defparam \_T_3557~5 .lut_mask = 16'h8008;
defparam \_T_3557~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3557~6 (
	.dataa(\ex_ctrl_mem_wr.01~q ),
	.datab(\_T_3557~2_combout ),
	.datac(\_T_3557~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\_T_3557~6_combout ),
	.cout());
defparam \_T_3557~6 .lut_mask = 16'hA8A8;
defparam \_T_3557~6 .sum_lutc_input = "datac";

dffeas \ex_csr_cmd[2] (
	.clk(clk_clk),
	.d(\ex_ctrl_csr_cmd~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_cmd[2]~q ),
	.prn(vcc));
defparam \ex_csr_cmd[2] .is_wysiwyg = "true";
defparam \ex_csr_cmd[2] .power_up = "low";

dffeas \ex_csr_cmd[0] (
	.clk(clk_clk),
	.d(\ex_csr_cmd~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_cmd[0]~q ),
	.prn(vcc));
defparam \ex_csr_cmd[0] .is_wysiwyg = "true";
defparam \ex_csr_cmd[0] .power_up = "low";

dffeas \ex_csr_cmd[1] (
	.clk(clk_clk),
	.d(\ex_csr_cmd~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_cmd[1]~q ),
	.prn(vcc));
defparam \ex_csr_cmd[1] .is_wysiwyg = "true";
defparam \ex_csr_cmd[1] .power_up = "low";

cyclone10lp_lcell_comb \alu_io_op1[23]~60 (
	.dataa(\ex_pc[23]~q ),
	.datab(\ex_reg_rs1_bypass[23]~121_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[23]~60_combout ),
	.cout());
defparam \alu_io_op1[23]~60 .lut_mask = 16'hAACC;
defparam \alu_io_op1[23]~60 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[27]~61 (
	.dataa(\ex_pc[27]~q ),
	.datab(\ex_reg_rs1_bypass[27]~137_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[27]~61_combout ),
	.cout());
defparam \alu_io_op1[27]~61 .lut_mask = 16'hAACC;
defparam \alu_io_op1[27]~61 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_legal~2 (
	.dataa(\Equal51~0_combout ),
	.datab(\ex_ctrl_legal~3_combout ),
	.datac(\ex_ctrl_mask_type~0_combout ),
	.datad(\ex_ctrl_csr_cmd~13_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_legal~2_combout ),
	.cout());
defparam \ex_ctrl_legal~2 .lut_mask = 16'hEFFF;
defparam \ex_ctrl_legal~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_GEN_32~0 (
	.dataa(\id_inst[12]~q ),
	.datab(gnd),
	.datac(\Equal11~0_combout ),
	.datad(\id_ctrl_br_type[2]~5_combout ),
	.cin(gnd),
	.combout(\_GEN_32~0_combout ),
	.cout());
defparam \_GEN_32~0 .lut_mask = 16'h00AF;
defparam \_GEN_32~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_GEN_32~1 (
	.dataa(\_T_1778~combout ),
	.datab(\_GEN_32~0_combout ),
	.datac(\id_ctrl_br_type[0]~9_combout ),
	.datad(\id_ctrl_br_type[1]~10_combout ),
	.cin(gnd),
	.combout(\_GEN_32~1_combout ),
	.cout());
defparam \_GEN_32~1 .lut_mask = 16'h0880;
defparam \_GEN_32~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[31]~62 (
	.dataa(\ex_pc[31]~q ),
	.datab(\ex_reg_rs1_bypass[31]~33_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[31]~62_combout ),
	.cout());
defparam \alu_io_op1[31]~62 .lut_mask = 16'hAACC;
defparam \alu_io_op1[31]~62 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_alu_op1[0]~5 (
	.dataa(\ex_reg_rs1_bypass[0]~16_combout ),
	.datab(\ex_npc[0]~q ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[0]~q ),
	.cin(gnd),
	.combout(\csr_io_alu_op1[0]~5_combout ),
	.cout());
defparam \csr_io_alu_op1[0]~5 .lut_mask = 16'hAACC;
defparam \csr_io_alu_op1[0]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[30]~63 (
	.dataa(\ex_pc[30]~q ),
	.datab(\ex_reg_rs1_bypass[30]~29_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[30]~63_combout ),
	.cout());
defparam \alu_io_op1[30]~63 .lut_mask = 16'hAACC;
defparam \alu_io_op1[30]~63 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_alu_op1[1]~6 (
	.dataa(\ex_reg_rs1_bypass[1]~11_combout ),
	.datab(\ex_npc[1]~q ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[0]~q ),
	.cin(gnd),
	.combout(\csr_io_alu_op1[1]~6_combout ),
	.cout());
defparam \csr_io_alu_op1[1]~6 .lut_mask = 16'hAACC;
defparam \csr_io_alu_op1[1]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[8]~64 (
	.dataa(\ex_pc[8]~q ),
	.datab(\ex_reg_rs1_bypass[8]~37_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[8]~64_combout ),
	.cout());
defparam \alu_io_op1[8]~64 .lut_mask = 16'hAACC;
defparam \alu_io_op1[8]~64 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[7]~65 (
	.dataa(\ex_pc[7]~q ),
	.datab(\ex_reg_rs1_bypass[7]~105_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[7]~65_combout ),
	.cout());
defparam \alu_io_op1[7]~65 .lut_mask = 16'hAACC;
defparam \alu_io_op1[7]~65 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[24]~66 (
	.dataa(\ex_pc[24]~q ),
	.datab(\ex_reg_rs1_bypass[24]~125_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[24]~66_combout ),
	.cout());
defparam \alu_io_op1[24]~66 .lut_mask = 16'hAACC;
defparam \alu_io_op1[24]~66 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[4]~67 (
	.dataa(\ex_pc[4]~q ),
	.datab(\ex_reg_rs1_bypass[4]~85_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[4]~67_combout ),
	.cout());
defparam \alu_io_op1[4]~67 .lut_mask = 16'hAACC;
defparam \alu_io_op1[4]~67 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[3]~68 (
	.dataa(\ex_pc[3]~q ),
	.datab(\ex_reg_rs1_bypass[3]~97_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[3]~68_combout ),
	.cout());
defparam \alu_io_op1[3]~68 .lut_mask = 16'hAACC;
defparam \alu_io_op1[3]~68 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[28]~69 (
	.dataa(\ex_pc[28]~q ),
	.datab(\ex_reg_rs1_bypass[28]~21_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[28]~69_combout ),
	.cout());
defparam \alu_io_op1[28]~69 .lut_mask = 16'hAACC;
defparam \alu_io_op1[28]~69 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[6]~70 (
	.dataa(\ex_pc[6]~q ),
	.datab(\ex_reg_rs1_bypass[6]~101_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[6]~70_combout ),
	.cout());
defparam \alu_io_op1[6]~70 .lut_mask = 16'hAACC;
defparam \alu_io_op1[6]~70 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[25]~71 (
	.dataa(\ex_pc[25]~q ),
	.datab(\ex_reg_rs1_bypass[25]~129_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[25]~71_combout ),
	.cout());
defparam \alu_io_op1[25]~71 .lut_mask = 16'hAACC;
defparam \alu_io_op1[25]~71 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[5]~72 (
	.dataa(\ex_pc[5]~q ),
	.datab(\ex_reg_rs1_bypass[5]~93_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[5]~72_combout ),
	.cout());
defparam \alu_io_op1[5]~72 .lut_mask = 16'hAACC;
defparam \alu_io_op1[5]~72 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[26]~73 (
	.dataa(\ex_pc[26]~q ),
	.datab(\ex_reg_rs1_bypass[26]~133_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[26]~73_combout ),
	.cout());
defparam \alu_io_op1[26]~73 .lut_mask = 16'hAACC;
defparam \alu_io_op1[26]~73 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[2]~74 (
	.dataa(\ex_pc[2]~q ),
	.datab(\ex_reg_rs1_bypass[2]~89_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[2]~74_combout ),
	.cout());
defparam \alu_io_op1[2]~74 .lut_mask = 16'hAACC;
defparam \alu_io_op1[2]~74 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[29]~75 (
	.dataa(\ex_pc[29]~q ),
	.datab(\ex_reg_rs1_bypass[29]~25_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[29]~75_combout ),
	.cout());
defparam \alu_io_op1[29]~75 .lut_mask = 16'hAACC;
defparam \alu_io_op1[29]~75 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[12]~76 (
	.dataa(\ex_pc[12]~q ),
	.datab(\ex_reg_rs1_bypass[12]~53_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[12]~76_combout ),
	.cout());
defparam \alu_io_op1[12]~76 .lut_mask = 16'hAACC;
defparam \alu_io_op1[12]~76 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[19]~77 (
	.dataa(\ex_pc[19]~q ),
	.datab(\ex_reg_rs1_bypass[19]~81_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[19]~77_combout ),
	.cout());
defparam \alu_io_op1[19]~77 .lut_mask = 16'hAACC;
defparam \alu_io_op1[19]~77 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[11]~78 (
	.dataa(\ex_pc[11]~q ),
	.datab(\ex_reg_rs1_bypass[11]~49_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[11]~78_combout ),
	.cout());
defparam \alu_io_op1[11]~78 .lut_mask = 16'hAACC;
defparam \alu_io_op1[11]~78 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[20]~79 (
	.dataa(\ex_pc[20]~q ),
	.datab(\ex_reg_rs1_bypass[20]~109_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[20]~79_combout ),
	.cout());
defparam \alu_io_op1[20]~79 .lut_mask = 16'hAACC;
defparam \alu_io_op1[20]~79 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[10]~80 (
	.dataa(\ex_pc[10]~q ),
	.datab(\ex_reg_rs1_bypass[10]~45_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[10]~80_combout ),
	.cout());
defparam \alu_io_op1[10]~80 .lut_mask = 16'hAACC;
defparam \alu_io_op1[10]~80 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[21]~81 (
	.dataa(\ex_pc[21]~q ),
	.datab(\ex_reg_rs1_bypass[21]~113_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[21]~81_combout ),
	.cout());
defparam \alu_io_op1[21]~81 .lut_mask = 16'hAACC;
defparam \alu_io_op1[21]~81 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[9]~82 (
	.dataa(\ex_pc[9]~q ),
	.datab(\ex_reg_rs1_bypass[9]~41_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[9]~82_combout ),
	.cout());
defparam \alu_io_op1[9]~82 .lut_mask = 16'hAACC;
defparam \alu_io_op1[9]~82 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[22]~83 (
	.dataa(\ex_pc[22]~q ),
	.datab(\ex_reg_rs1_bypass[22]~117_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[22]~83_combout ),
	.cout());
defparam \alu_io_op1[22]~83 .lut_mask = 16'hAACC;
defparam \alu_io_op1[22]~83 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[16]~84 (
	.dataa(\ex_pc[16]~q ),
	.datab(\ex_reg_rs1_bypass[16]~69_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[16]~84_combout ),
	.cout());
defparam \alu_io_op1[16]~84 .lut_mask = 16'hAACC;
defparam \alu_io_op1[16]~84 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[15]~85 (
	.dataa(\ex_pc[15]~q ),
	.datab(\ex_reg_rs1_bypass[15]~65_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[15]~85_combout ),
	.cout());
defparam \alu_io_op1[15]~85 .lut_mask = 16'hAACC;
defparam \alu_io_op1[15]~85 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[14]~86 (
	.dataa(\ex_pc[14]~q ),
	.datab(\ex_reg_rs1_bypass[14]~61_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[14]~86_combout ),
	.cout());
defparam \alu_io_op1[14]~86 .lut_mask = 16'hAACC;
defparam \alu_io_op1[14]~86 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[17]~87 (
	.dataa(\ex_pc[17]~q ),
	.datab(\ex_reg_rs1_bypass[17]~73_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[17]~87_combout ),
	.cout());
defparam \alu_io_op1[17]~87 .lut_mask = 16'hAACC;
defparam \alu_io_op1[17]~87 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[13]~88 (
	.dataa(\ex_pc[13]~q ),
	.datab(\ex_reg_rs1_bypass[13]~57_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[13]~88_combout ),
	.cout());
defparam \alu_io_op1[13]~88 .lut_mask = 16'hAACC;
defparam \alu_io_op1[13]~88 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[18]~89 (
	.dataa(\ex_pc[18]~q ),
	.datab(\ex_reg_rs1_bypass[18]~77_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_op1[1]~q ),
	.cin(gnd),
	.combout(\alu_io_op1[18]~89_combout ),
	.cout());
defparam \alu_io_op1[18]~89 .lut_mask = 16'hAACC;
defparam \alu_io_op1[18]~89 .sum_lutc_input = "datac";

dffeas wb_dmem_read_ack(
	.clk(clk_clk),
	.d(\wb_dmem_read_ack~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_ack~q ),
	.prn(vcc));
defparam wb_dmem_read_ack.is_wysiwyg = "true";
defparam wb_dmem_read_ack.power_up = "low";

cyclone10lp_lcell_comb _GEN_9(
	.dataa(mem_ctrl_mem_wr01),
	.datab(\_T_3549~q ),
	.datac(gnd),
	.datad(\wb_dmem_read_ack~q ),
	.cin(gnd),
	.combout(\_GEN_9~combout ),
	.cout());
defparam _GEN_9.lut_mask = 16'hAAEE;
defparam _GEN_9.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_csr_cmd~15 (
	.dataa(\ex_ctrl_mask_type~0_combout ),
	.datab(\Equal51~0_combout ),
	.datac(\ex_ctrl_wb_sel~12_combout ),
	.datad(\ex_ctrl_csr_cmd~13_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_csr_cmd~15_combout ),
	.cout());
defparam \ex_ctrl_csr_cmd~15 .lut_mask = 16'h88A0;
defparam \ex_ctrl_csr_cmd~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal47~0 (
	.dataa(\id_inst[4]~q ),
	.datab(\id_inst[6]~q ),
	.datac(\id_inst[12]~q ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\Equal47~0_combout ),
	.cout());
defparam \Equal47~0 .lut_mask = 16'h8000;
defparam \Equal47~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_csr_cmd~6 (
	.dataa(\ex_ctrl_csr_cmd~9_combout ),
	.datab(\ex_ctrl_csr_cmd~11_combout ),
	.datac(\Equal13~0_combout ),
	.datad(\Equal43~0_combout ),
	.cin(gnd),
	.combout(\ex_csr_cmd~6_combout ),
	.cout());
defparam \ex_csr_cmd~6 .lut_mask = 16'h0888;
defparam \ex_csr_cmd~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_csr_cmd~7 (
	.dataa(\ex_ctrl_mask_type~0_combout ),
	.datab(\Equal47~0_combout ),
	.datac(\ex_csr_cmd~6_combout ),
	.datad(\ex_ctrl_csr_cmd~12_combout ),
	.cin(gnd),
	.combout(\ex_csr_cmd~7_combout ),
	.cout());
defparam \ex_csr_cmd~7 .lut_mask = 16'h88A0;
defparam \ex_csr_cmd~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_csr_cmd~8 (
	.dataa(\id_inst[13]~q ),
	.datab(\Equal43~0_combout ),
	.datac(\ex_csr_cmd~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_csr_cmd~8_combout ),
	.cout());
defparam \ex_csr_cmd~8 .lut_mask = 16'h8080;
defparam \ex_csr_cmd~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_csr_cmd~9 (
	.dataa(\ex_ctrl_mask_type~0_combout ),
	.datab(\ex_csr_cmd~8_combout ),
	.datac(\ex_ctrl_csr_cmd~12_combout ),
	.datad(\ex_csr_cmd~4_combout ),
	.cin(gnd),
	.combout(\ex_csr_cmd~9_combout ),
	.cout());
defparam \ex_csr_cmd~9 .lut_mask = 16'h08A8;
defparam \ex_csr_cmd~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_sw_r_ex_imm[0]~9 (
	.dataa(\ex_inst[7]~q ),
	.datab(\io_sw_r_ex_imm[0]~2_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_imm_type.001~q ),
	.cin(gnd),
	.combout(\io_sw_r_ex_imm[0]~9_combout ),
	.cout());
defparam \io_sw_r_ex_imm[0]~9 .lut_mask = 16'hAACC;
defparam \io_sw_r_ex_imm[0]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[0]~1 (
	.dataa(\Equal60~5_combout ),
	.datab(\wb_ctrl_csr_cmd.000~q ),
	.datac(\Equal61~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_io_in[0]~1_combout ),
	.cout());
defparam \csr_io_in[0]~1 .lut_mask = 16'hEAEA;
defparam \csr_io_in[0]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[0]~2 (
	.dataa(\Equal61~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal60~5_combout ),
	.cin(gnd),
	.combout(\csr_io_in[0]~2_combout ),
	.cout());
defparam \csr_io_in[0]~2 .lut_mask = 16'h00AA;
defparam \csr_io_in[0]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[0]~3 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[0]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[0]~16_combout ),
	.cin(gnd),
	.combout(\csr_io_in[0]~3_combout ),
	.cout());
defparam \csr_io_in[0]~3 .lut_mask = 16'hE5E0;
defparam \csr_io_in[0]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[0]~4 (
	.dataa(mem_alu_out_0),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[0]~3_combout ),
	.datad(\wb_csr_data[0]~q ),
	.cin(gnd),
	.combout(\csr_io_in[0]~4_combout ),
	.cout());
defparam \csr_io_in[0]~4 .lut_mask = 16'hF838;
defparam \csr_io_in[0]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[0]~5 (
	.dataa(\mem_csr_data[0]~q ),
	.datab(\csr_io_in[0]~4_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[0]~5_combout ),
	.cout());
defparam \csr_io_in[0]~5 .lut_mask = 16'h00AC;
defparam \csr_io_in[0]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[0]~6 (
	.dataa(\csr_io_in[0]~5_combout ),
	.datab(\ex_ctrl_imm_type.101~q ),
	.datac(\io_sw_r_ex_imm[0]~9_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_io_in[0]~6_combout ),
	.cout());
defparam \csr_io_in[0]~6 .lut_mask = 16'hEAEA;
defparam \csr_io_in[0]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[1]~7 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(mem_alu_out_1),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[1]~11_combout ),
	.cin(gnd),
	.combout(\csr_io_in[1]~7_combout ),
	.cout());
defparam \csr_io_in[1]~7 .lut_mask = 16'hE5E0;
defparam \csr_io_in[1]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[1]~8 (
	.dataa(\wb_alu_out[1]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[1]~7_combout ),
	.datad(\wb_csr_data[1]~q ),
	.cin(gnd),
	.combout(\csr_io_in[1]~8_combout ),
	.cout());
defparam \csr_io_in[1]~8 .lut_mask = 16'hF838;
defparam \csr_io_in[1]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[1]~9 (
	.dataa(\mem_csr_data[1]~q ),
	.datab(\csr_io_in[1]~8_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[1]~9_combout ),
	.cout());
defparam \csr_io_in[1]~9 .lut_mask = 16'h00AC;
defparam \csr_io_in[1]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[1]~10 (
	.dataa(\csr_io_in[1]~9_combout ),
	.datab(\ex_ctrl_imm_type.101~q ),
	.datac(\io_sw_r_ex_imm[1]~1_combout ),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\csr_io_in[1]~10_combout ),
	.cout());
defparam \csr_io_in[1]~10 .lut_mask = 16'hAAEA;
defparam \csr_io_in[1]~10 .sum_lutc_input = "datac";

dffeas \ex_inst[0] (
	.clk(clk_clk),
	.d(\ex_inst~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[0]~q ),
	.prn(vcc));
defparam \ex_inst[0] .is_wysiwyg = "true";
defparam \ex_inst[0] .power_up = "low";

dffeas \ex_inst[1] (
	.clk(clk_clk),
	.d(\ex_inst~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[1]~q ),
	.prn(vcc));
defparam \ex_inst[1] .is_wysiwyg = "true";
defparam \ex_inst[1] .power_up = "low";

dffeas \ex_inst[4] (
	.clk(clk_clk),
	.d(\ex_inst~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[4]~q ),
	.prn(vcc));
defparam \ex_inst[4] .is_wysiwyg = "true";
defparam \ex_inst[4] .power_up = "low";

dffeas \ex_inst[2] (
	.clk(clk_clk),
	.d(\ex_inst~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[2]~q ),
	.prn(vcc));
defparam \ex_inst[2] .is_wysiwyg = "true";
defparam \ex_inst[2] .power_up = "low";

dffeas \ex_inst[3] (
	.clk(clk_clk),
	.d(\ex_inst~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[3]~q ),
	.prn(vcc));
defparam \ex_inst[3] .is_wysiwyg = "true";
defparam \ex_inst[3] .power_up = "low";

dffeas \ex_inst[5] (
	.clk(clk_clk),
	.d(\ex_inst~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[5]~q ),
	.prn(vcc));
defparam \ex_inst[5] .is_wysiwyg = "true";
defparam \ex_inst[5] .power_up = "low";

dffeas \ex_inst[6] (
	.clk(clk_clk),
	.d(\ex_inst~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[6]~q ),
	.prn(vcc));
defparam \ex_inst[6] .is_wysiwyg = "true";
defparam \ex_inst[6] .power_up = "low";

cyclone10lp_lcell_comb \wb_dmem_read_ack~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(read_latency_shift_reg_01),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_dmem_read_ack~0_combout ),
	.cout());
defparam \wb_dmem_read_ack~0 .lut_mask = 16'h8888;
defparam \wb_dmem_read_ack~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[2]~11 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[2]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[2]~89_combout ),
	.cin(gnd),
	.combout(\csr_io_in[2]~11_combout ),
	.cout());
defparam \csr_io_in[2]~11 .lut_mask = 16'hE5E0;
defparam \csr_io_in[2]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[2]~12 (
	.dataa(mem_alu_out_2),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[2]~11_combout ),
	.datad(\wb_csr_data[2]~q ),
	.cin(gnd),
	.combout(\csr_io_in[2]~12_combout ),
	.cout());
defparam \csr_io_in[2]~12 .lut_mask = 16'hF838;
defparam \csr_io_in[2]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[2]~13 (
	.dataa(\mem_csr_data[2]~q ),
	.datab(\csr_io_in[2]~12_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[2]~13_combout ),
	.cout());
defparam \csr_io_in[2]~13 .lut_mask = 16'h00AC;
defparam \csr_io_in[2]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[2]~14 (
	.dataa(\csr_io_in[2]~13_combout ),
	.datab(\ex_ctrl_imm_type.101~q ),
	.datac(\io_sw_r_ex_imm[2]~6_combout ),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\csr_io_in[2]~14_combout ),
	.cout());
defparam \csr_io_in[2]~14 .lut_mask = 16'hAAEA;
defparam \csr_io_in[2]~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[3]~15 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(mem_alu_out_3),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[3]~97_combout ),
	.cin(gnd),
	.combout(\csr_io_in[3]~15_combout ),
	.cout());
defparam \csr_io_in[3]~15 .lut_mask = 16'hE5E0;
defparam \csr_io_in[3]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[3]~16 (
	.dataa(\wb_alu_out[3]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[3]~15_combout ),
	.datad(\wb_csr_data[3]~q ),
	.cin(gnd),
	.combout(\csr_io_in[3]~16_combout ),
	.cout());
defparam \csr_io_in[3]~16 .lut_mask = 16'hF838;
defparam \csr_io_in[3]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[3]~17 (
	.dataa(\mem_csr_data[3]~q ),
	.datab(\csr_io_in[3]~16_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[3]~17_combout ),
	.cout());
defparam \csr_io_in[3]~17 .lut_mask = 16'h00AC;
defparam \csr_io_in[3]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[3]~18 (
	.dataa(\csr_io_in[3]~17_combout ),
	.datab(\ex_ctrl_imm_type.101~q ),
	.datac(\io_sw_r_ex_imm[3]~8_combout ),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\csr_io_in[3]~18_combout ),
	.cout());
defparam \csr_io_in[3]~18 .lut_mask = 16'hAAEA;
defparam \csr_io_in[3]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[4]~19 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[4]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[4]~85_combout ),
	.cin(gnd),
	.combout(\csr_io_in[4]~19_combout ),
	.cout());
defparam \csr_io_in[4]~19 .lut_mask = 16'hE5E0;
defparam \csr_io_in[4]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[4]~20 (
	.dataa(\mem_alu_out[4]~q ),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[4]~19_combout ),
	.datad(\wb_csr_data[4]~q ),
	.cin(gnd),
	.combout(\csr_io_in[4]~20_combout ),
	.cout());
defparam \csr_io_in[4]~20 .lut_mask = 16'hF838;
defparam \csr_io_in[4]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[4]~21 (
	.dataa(\mem_csr_data[4]~q ),
	.datab(\csr_io_in[4]~20_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[4]~21_combout ),
	.cout());
defparam \csr_io_in[4]~21 .lut_mask = 16'h00AC;
defparam \csr_io_in[4]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[4]~22 (
	.dataa(\csr_io_in[4]~21_combout ),
	.datab(\ex_ctrl_imm_type.101~q ),
	.datac(\io_sw_r_ex_imm[4]~4_combout ),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\csr_io_in[4]~22_combout ),
	.cout());
defparam \csr_io_in[4]~22 .lut_mask = 16'hAAEA;
defparam \csr_io_in[4]~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[5]~23 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(\mem_alu_out[5]~q ),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[5]~93_combout ),
	.cin(gnd),
	.combout(\csr_io_in[5]~23_combout ),
	.cout());
defparam \csr_io_in[5]~23 .lut_mask = 16'hE5E0;
defparam \csr_io_in[5]~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[5]~24 (
	.dataa(\wb_alu_out[5]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[5]~23_combout ),
	.datad(\wb_csr_data[5]~q ),
	.cin(gnd),
	.combout(\csr_io_in[5]~24_combout ),
	.cout());
defparam \csr_io_in[5]~24 .lut_mask = 16'hF838;
defparam \csr_io_in[5]~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[5]~25 (
	.dataa(\mem_csr_data[5]~q ),
	.datab(\csr_io_in[5]~24_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[5]~25_combout ),
	.cout());
defparam \csr_io_in[5]~25 .lut_mask = 16'h00AC;
defparam \csr_io_in[5]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[6]~26 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[6]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[6]~101_combout ),
	.cin(gnd),
	.combout(\csr_io_in[6]~26_combout ),
	.cout());
defparam \csr_io_in[6]~26 .lut_mask = 16'hE5E0;
defparam \csr_io_in[6]~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[6]~27 (
	.dataa(\mem_alu_out[6]~q ),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[6]~26_combout ),
	.datad(\wb_csr_data[6]~q ),
	.cin(gnd),
	.combout(\csr_io_in[6]~27_combout ),
	.cout());
defparam \csr_io_in[6]~27 .lut_mask = 16'hF838;
defparam \csr_io_in[6]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[6]~28 (
	.dataa(\mem_csr_data[6]~q ),
	.datab(\csr_io_in[6]~27_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[6]~28_combout ),
	.cout());
defparam \csr_io_in[6]~28 .lut_mask = 16'h00AC;
defparam \csr_io_in[6]~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[7]~29 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(\mem_alu_out[7]~q ),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[7]~105_combout ),
	.cin(gnd),
	.combout(\csr_io_in[7]~29_combout ),
	.cout());
defparam \csr_io_in[7]~29 .lut_mask = 16'hE5E0;
defparam \csr_io_in[7]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[7]~30 (
	.dataa(\wb_alu_out[7]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[7]~29_combout ),
	.datad(\wb_csr_data[7]~q ),
	.cin(gnd),
	.combout(\csr_io_in[7]~30_combout ),
	.cout());
defparam \csr_io_in[7]~30 .lut_mask = 16'hF838;
defparam \csr_io_in[7]~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[7]~31 (
	.dataa(\mem_csr_data[7]~q ),
	.datab(\csr_io_in[7]~30_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[7]~31_combout ),
	.cout());
defparam \csr_io_in[7]~31 .lut_mask = 16'h00AC;
defparam \csr_io_in[7]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[8]~32 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[8]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[8]~37_combout ),
	.cin(gnd),
	.combout(\csr_io_in[8]~32_combout ),
	.cout());
defparam \csr_io_in[8]~32 .lut_mask = 16'hE5E0;
defparam \csr_io_in[8]~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[8]~33 (
	.dataa(\mem_alu_out[8]~q ),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[8]~32_combout ),
	.datad(\wb_csr_data[8]~q ),
	.cin(gnd),
	.combout(\csr_io_in[8]~33_combout ),
	.cout());
defparam \csr_io_in[8]~33 .lut_mask = 16'hF838;
defparam \csr_io_in[8]~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[8]~34 (
	.dataa(\mem_csr_data[8]~q ),
	.datab(\csr_io_in[8]~33_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[8]~34_combout ),
	.cout());
defparam \csr_io_in[8]~34 .lut_mask = 16'h00AC;
defparam \csr_io_in[8]~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[9]~35 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(\mem_alu_out[9]~q ),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[9]~41_combout ),
	.cin(gnd),
	.combout(\csr_io_in[9]~35_combout ),
	.cout());
defparam \csr_io_in[9]~35 .lut_mask = 16'hE5E0;
defparam \csr_io_in[9]~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[9]~36 (
	.dataa(\wb_alu_out[9]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[9]~35_combout ),
	.datad(\wb_csr_data[9]~q ),
	.cin(gnd),
	.combout(\csr_io_in[9]~36_combout ),
	.cout());
defparam \csr_io_in[9]~36 .lut_mask = 16'hF838;
defparam \csr_io_in[9]~36 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[9]~37 (
	.dataa(\mem_csr_data[9]~q ),
	.datab(\csr_io_in[9]~36_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[9]~37_combout ),
	.cout());
defparam \csr_io_in[9]~37 .lut_mask = 16'h00AC;
defparam \csr_io_in[9]~37 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[10]~38 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[10]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[10]~45_combout ),
	.cin(gnd),
	.combout(\csr_io_in[10]~38_combout ),
	.cout());
defparam \csr_io_in[10]~38 .lut_mask = 16'hE5E0;
defparam \csr_io_in[10]~38 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[10]~39 (
	.dataa(\mem_alu_out[10]~q ),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[10]~38_combout ),
	.datad(\wb_csr_data[10]~q ),
	.cin(gnd),
	.combout(\csr_io_in[10]~39_combout ),
	.cout());
defparam \csr_io_in[10]~39 .lut_mask = 16'hF838;
defparam \csr_io_in[10]~39 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[10]~40 (
	.dataa(\mem_csr_data[10]~q ),
	.datab(\csr_io_in[10]~39_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[10]~40_combout ),
	.cout());
defparam \csr_io_in[10]~40 .lut_mask = 16'h00AC;
defparam \csr_io_in[10]~40 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[11]~41 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(\mem_alu_out[11]~q ),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[11]~49_combout ),
	.cin(gnd),
	.combout(\csr_io_in[11]~41_combout ),
	.cout());
defparam \csr_io_in[11]~41 .lut_mask = 16'hE5E0;
defparam \csr_io_in[11]~41 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[11]~42 (
	.dataa(\wb_alu_out[11]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[11]~41_combout ),
	.datad(\wb_csr_data[11]~q ),
	.cin(gnd),
	.combout(\csr_io_in[11]~42_combout ),
	.cout());
defparam \csr_io_in[11]~42 .lut_mask = 16'hF838;
defparam \csr_io_in[11]~42 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[11]~43 (
	.dataa(\mem_csr_data[11]~q ),
	.datab(\csr_io_in[11]~42_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[11]~43_combout ),
	.cout());
defparam \csr_io_in[11]~43 .lut_mask = 16'h00AC;
defparam \csr_io_in[11]~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[12]~44 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[12]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[12]~53_combout ),
	.cin(gnd),
	.combout(\csr_io_in[12]~44_combout ),
	.cout());
defparam \csr_io_in[12]~44 .lut_mask = 16'hE5E0;
defparam \csr_io_in[12]~44 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[12]~45 (
	.dataa(\mem_alu_out[12]~q ),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[12]~44_combout ),
	.datad(\wb_csr_data[12]~q ),
	.cin(gnd),
	.combout(\csr_io_in[12]~45_combout ),
	.cout());
defparam \csr_io_in[12]~45 .lut_mask = 16'hF838;
defparam \csr_io_in[12]~45 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[12]~46 (
	.dataa(\mem_csr_data[12]~q ),
	.datab(\csr_io_in[12]~45_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[12]~46_combout ),
	.cout());
defparam \csr_io_in[12]~46 .lut_mask = 16'h00AC;
defparam \csr_io_in[12]~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[13]~47 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(\mem_alu_out[13]~q ),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[13]~57_combout ),
	.cin(gnd),
	.combout(\csr_io_in[13]~47_combout ),
	.cout());
defparam \csr_io_in[13]~47 .lut_mask = 16'hE5E0;
defparam \csr_io_in[13]~47 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[13]~48 (
	.dataa(\wb_alu_out[13]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[13]~47_combout ),
	.datad(\wb_csr_data[13]~q ),
	.cin(gnd),
	.combout(\csr_io_in[13]~48_combout ),
	.cout());
defparam \csr_io_in[13]~48 .lut_mask = 16'hF838;
defparam \csr_io_in[13]~48 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[13]~49 (
	.dataa(\mem_csr_data[13]~q ),
	.datab(\csr_io_in[13]~48_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[13]~49_combout ),
	.cout());
defparam \csr_io_in[13]~49 .lut_mask = 16'h00AC;
defparam \csr_io_in[13]~49 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[14]~50 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[14]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[14]~61_combout ),
	.cin(gnd),
	.combout(\csr_io_in[14]~50_combout ),
	.cout());
defparam \csr_io_in[14]~50 .lut_mask = 16'hE5E0;
defparam \csr_io_in[14]~50 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[14]~51 (
	.dataa(\mem_alu_out[14]~q ),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[14]~50_combout ),
	.datad(\wb_csr_data[14]~q ),
	.cin(gnd),
	.combout(\csr_io_in[14]~51_combout ),
	.cout());
defparam \csr_io_in[14]~51 .lut_mask = 16'hF838;
defparam \csr_io_in[14]~51 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[14]~52 (
	.dataa(\mem_csr_data[14]~q ),
	.datab(\csr_io_in[14]~51_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[14]~52_combout ),
	.cout());
defparam \csr_io_in[14]~52 .lut_mask = 16'h00AC;
defparam \csr_io_in[14]~52 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[15]~53 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(\mem_alu_out[15]~q ),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[15]~65_combout ),
	.cin(gnd),
	.combout(\csr_io_in[15]~53_combout ),
	.cout());
defparam \csr_io_in[15]~53 .lut_mask = 16'hE5E0;
defparam \csr_io_in[15]~53 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[15]~54 (
	.dataa(\wb_alu_out[15]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[15]~53_combout ),
	.datad(\wb_csr_data[15]~q ),
	.cin(gnd),
	.combout(\csr_io_in[15]~54_combout ),
	.cout());
defparam \csr_io_in[15]~54 .lut_mask = 16'hF838;
defparam \csr_io_in[15]~54 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[15]~55 (
	.dataa(\mem_csr_data[15]~q ),
	.datab(\csr_io_in[15]~54_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[15]~55_combout ),
	.cout());
defparam \csr_io_in[15]~55 .lut_mask = 16'h00AC;
defparam \csr_io_in[15]~55 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[16]~56 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[16]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[16]~69_combout ),
	.cin(gnd),
	.combout(\csr_io_in[16]~56_combout ),
	.cout());
defparam \csr_io_in[16]~56 .lut_mask = 16'hE5E0;
defparam \csr_io_in[16]~56 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[16]~57 (
	.dataa(\mem_alu_out[16]~q ),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[16]~56_combout ),
	.datad(\wb_csr_data[16]~q ),
	.cin(gnd),
	.combout(\csr_io_in[16]~57_combout ),
	.cout());
defparam \csr_io_in[16]~57 .lut_mask = 16'hF838;
defparam \csr_io_in[16]~57 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[16]~58 (
	.dataa(\mem_csr_data[16]~q ),
	.datab(\csr_io_in[16]~57_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[16]~58_combout ),
	.cout());
defparam \csr_io_in[16]~58 .lut_mask = 16'h00AC;
defparam \csr_io_in[16]~58 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[17]~59 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(\mem_alu_out[17]~q ),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[17]~73_combout ),
	.cin(gnd),
	.combout(\csr_io_in[17]~59_combout ),
	.cout());
defparam \csr_io_in[17]~59 .lut_mask = 16'hE5E0;
defparam \csr_io_in[17]~59 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[17]~60 (
	.dataa(\wb_alu_out[17]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[17]~59_combout ),
	.datad(\wb_csr_data[17]~q ),
	.cin(gnd),
	.combout(\csr_io_in[17]~60_combout ),
	.cout());
defparam \csr_io_in[17]~60 .lut_mask = 16'hF838;
defparam \csr_io_in[17]~60 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[17]~61 (
	.dataa(\mem_csr_data[17]~q ),
	.datab(\csr_io_in[17]~60_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[17]~61_combout ),
	.cout());
defparam \csr_io_in[17]~61 .lut_mask = 16'h00AC;
defparam \csr_io_in[17]~61 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[18]~62 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[18]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[18]~77_combout ),
	.cin(gnd),
	.combout(\csr_io_in[18]~62_combout ),
	.cout());
defparam \csr_io_in[18]~62 .lut_mask = 16'hE5E0;
defparam \csr_io_in[18]~62 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[18]~63 (
	.dataa(\mem_alu_out[18]~q ),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[18]~62_combout ),
	.datad(\wb_csr_data[18]~q ),
	.cin(gnd),
	.combout(\csr_io_in[18]~63_combout ),
	.cout());
defparam \csr_io_in[18]~63 .lut_mask = 16'hF838;
defparam \csr_io_in[18]~63 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[18]~64 (
	.dataa(\mem_csr_data[18]~q ),
	.datab(\csr_io_in[18]~63_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[18]~64_combout ),
	.cout());
defparam \csr_io_in[18]~64 .lut_mask = 16'h00AC;
defparam \csr_io_in[18]~64 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[19]~65 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(\mem_alu_out[19]~q ),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[19]~81_combout ),
	.cin(gnd),
	.combout(\csr_io_in[19]~65_combout ),
	.cout());
defparam \csr_io_in[19]~65 .lut_mask = 16'hE5E0;
defparam \csr_io_in[19]~65 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[19]~66 (
	.dataa(\wb_alu_out[19]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[19]~65_combout ),
	.datad(\wb_csr_data[19]~q ),
	.cin(gnd),
	.combout(\csr_io_in[19]~66_combout ),
	.cout());
defparam \csr_io_in[19]~66 .lut_mask = 16'hF838;
defparam \csr_io_in[19]~66 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[19]~67 (
	.dataa(\mem_csr_data[19]~q ),
	.datab(\csr_io_in[19]~66_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[19]~67_combout ),
	.cout());
defparam \csr_io_in[19]~67 .lut_mask = 16'h00AC;
defparam \csr_io_in[19]~67 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[20]~68 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[20]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[20]~109_combout ),
	.cin(gnd),
	.combout(\csr_io_in[20]~68_combout ),
	.cout());
defparam \csr_io_in[20]~68 .lut_mask = 16'hE5E0;
defparam \csr_io_in[20]~68 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[20]~69 (
	.dataa(\mem_alu_out[20]~q ),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[20]~68_combout ),
	.datad(\wb_csr_data[20]~q ),
	.cin(gnd),
	.combout(\csr_io_in[20]~69_combout ),
	.cout());
defparam \csr_io_in[20]~69 .lut_mask = 16'hF838;
defparam \csr_io_in[20]~69 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[20]~70 (
	.dataa(\mem_csr_data[20]~q ),
	.datab(\csr_io_in[20]~69_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[20]~70_combout ),
	.cout());
defparam \csr_io_in[20]~70 .lut_mask = 16'h00AC;
defparam \csr_io_in[20]~70 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[21]~71 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(\mem_alu_out[21]~q ),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[21]~113_combout ),
	.cin(gnd),
	.combout(\csr_io_in[21]~71_combout ),
	.cout());
defparam \csr_io_in[21]~71 .lut_mask = 16'hE5E0;
defparam \csr_io_in[21]~71 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[21]~72 (
	.dataa(\wb_alu_out[21]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[21]~71_combout ),
	.datad(\wb_csr_data[21]~q ),
	.cin(gnd),
	.combout(\csr_io_in[21]~72_combout ),
	.cout());
defparam \csr_io_in[21]~72 .lut_mask = 16'hF838;
defparam \csr_io_in[21]~72 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[21]~73 (
	.dataa(\mem_csr_data[21]~q ),
	.datab(\csr_io_in[21]~72_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[21]~73_combout ),
	.cout());
defparam \csr_io_in[21]~73 .lut_mask = 16'h00AC;
defparam \csr_io_in[21]~73 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[22]~74 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[22]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[22]~117_combout ),
	.cin(gnd),
	.combout(\csr_io_in[22]~74_combout ),
	.cout());
defparam \csr_io_in[22]~74 .lut_mask = 16'hE5E0;
defparam \csr_io_in[22]~74 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[22]~75 (
	.dataa(\mem_alu_out[22]~q ),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[22]~74_combout ),
	.datad(\wb_csr_data[22]~q ),
	.cin(gnd),
	.combout(\csr_io_in[22]~75_combout ),
	.cout());
defparam \csr_io_in[22]~75 .lut_mask = 16'hF838;
defparam \csr_io_in[22]~75 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[22]~76 (
	.dataa(\mem_csr_data[22]~q ),
	.datab(\csr_io_in[22]~75_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[22]~76_combout ),
	.cout());
defparam \csr_io_in[22]~76 .lut_mask = 16'h00AC;
defparam \csr_io_in[22]~76 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[23]~77 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(\mem_alu_out[23]~q ),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[23]~121_combout ),
	.cin(gnd),
	.combout(\csr_io_in[23]~77_combout ),
	.cout());
defparam \csr_io_in[23]~77 .lut_mask = 16'hE5E0;
defparam \csr_io_in[23]~77 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[23]~78 (
	.dataa(\wb_alu_out[23]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[23]~77_combout ),
	.datad(\wb_csr_data[23]~q ),
	.cin(gnd),
	.combout(\csr_io_in[23]~78_combout ),
	.cout());
defparam \csr_io_in[23]~78 .lut_mask = 16'hF838;
defparam \csr_io_in[23]~78 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[23]~79 (
	.dataa(\mem_csr_data[23]~q ),
	.datab(\csr_io_in[23]~78_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[23]~79_combout ),
	.cout());
defparam \csr_io_in[23]~79 .lut_mask = 16'h00AC;
defparam \csr_io_in[23]~79 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[24]~80 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[24]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[24]~125_combout ),
	.cin(gnd),
	.combout(\csr_io_in[24]~80_combout ),
	.cout());
defparam \csr_io_in[24]~80 .lut_mask = 16'hE5E0;
defparam \csr_io_in[24]~80 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[24]~81 (
	.dataa(\mem_alu_out[24]~q ),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[24]~80_combout ),
	.datad(\wb_csr_data[24]~q ),
	.cin(gnd),
	.combout(\csr_io_in[24]~81_combout ),
	.cout());
defparam \csr_io_in[24]~81 .lut_mask = 16'hF838;
defparam \csr_io_in[24]~81 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[24]~82 (
	.dataa(\mem_csr_data[24]~q ),
	.datab(\csr_io_in[24]~81_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[24]~82_combout ),
	.cout());
defparam \csr_io_in[24]~82 .lut_mask = 16'h00AC;
defparam \csr_io_in[24]~82 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[25]~83 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(\mem_alu_out[25]~q ),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[25]~129_combout ),
	.cin(gnd),
	.combout(\csr_io_in[25]~83_combout ),
	.cout());
defparam \csr_io_in[25]~83 .lut_mask = 16'hE5E0;
defparam \csr_io_in[25]~83 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[25]~84 (
	.dataa(\wb_alu_out[25]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[25]~83_combout ),
	.datad(\wb_csr_data[25]~q ),
	.cin(gnd),
	.combout(\csr_io_in[25]~84_combout ),
	.cout());
defparam \csr_io_in[25]~84 .lut_mask = 16'hF838;
defparam \csr_io_in[25]~84 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[25]~85 (
	.dataa(\mem_csr_data[25]~q ),
	.datab(\csr_io_in[25]~84_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[25]~85_combout ),
	.cout());
defparam \csr_io_in[25]~85 .lut_mask = 16'h00AC;
defparam \csr_io_in[25]~85 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[26]~86 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[26]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[26]~133_combout ),
	.cin(gnd),
	.combout(\csr_io_in[26]~86_combout ),
	.cout());
defparam \csr_io_in[26]~86 .lut_mask = 16'hE5E0;
defparam \csr_io_in[26]~86 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[26]~87 (
	.dataa(\mem_alu_out[26]~q ),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[26]~86_combout ),
	.datad(\wb_csr_data[26]~q ),
	.cin(gnd),
	.combout(\csr_io_in[26]~87_combout ),
	.cout());
defparam \csr_io_in[26]~87 .lut_mask = 16'hF838;
defparam \csr_io_in[26]~87 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[26]~88 (
	.dataa(\mem_csr_data[26]~q ),
	.datab(\csr_io_in[26]~87_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[26]~88_combout ),
	.cout());
defparam \csr_io_in[26]~88 .lut_mask = 16'h00AC;
defparam \csr_io_in[26]~88 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[27]~89 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(\mem_alu_out[27]~q ),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[27]~137_combout ),
	.cin(gnd),
	.combout(\csr_io_in[27]~89_combout ),
	.cout());
defparam \csr_io_in[27]~89 .lut_mask = 16'hE5E0;
defparam \csr_io_in[27]~89 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[27]~90 (
	.dataa(\wb_alu_out[27]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[27]~89_combout ),
	.datad(\wb_csr_data[27]~q ),
	.cin(gnd),
	.combout(\csr_io_in[27]~90_combout ),
	.cout());
defparam \csr_io_in[27]~90 .lut_mask = 16'hF838;
defparam \csr_io_in[27]~90 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[27]~91 (
	.dataa(\mem_csr_data[27]~q ),
	.datab(\csr_io_in[27]~90_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[27]~91_combout ),
	.cout());
defparam \csr_io_in[27]~91 .lut_mask = 16'h00AC;
defparam \csr_io_in[27]~91 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[28]~92 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[28]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[28]~21_combout ),
	.cin(gnd),
	.combout(\csr_io_in[28]~92_combout ),
	.cout());
defparam \csr_io_in[28]~92 .lut_mask = 16'hE5E0;
defparam \csr_io_in[28]~92 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[28]~93 (
	.dataa(\mem_alu_out[28]~q ),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[28]~92_combout ),
	.datad(\wb_csr_data[28]~q ),
	.cin(gnd),
	.combout(\csr_io_in[28]~93_combout ),
	.cout());
defparam \csr_io_in[28]~93 .lut_mask = 16'hF838;
defparam \csr_io_in[28]~93 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[28]~94 (
	.dataa(\mem_csr_data[28]~q ),
	.datab(\csr_io_in[28]~93_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[28]~94_combout ),
	.cout());
defparam \csr_io_in[28]~94 .lut_mask = 16'h00AC;
defparam \csr_io_in[28]~94 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[29]~95 (
	.dataa(\csr_io_in[0]~2_combout ),
	.datab(\mem_alu_out[29]~q ),
	.datac(\csr_io_in[0]~1_combout ),
	.datad(\ex_reg_rs1_bypass[29]~25_combout ),
	.cin(gnd),
	.combout(\csr_io_in[29]~95_combout ),
	.cout());
defparam \csr_io_in[29]~95 .lut_mask = 16'hE5E0;
defparam \csr_io_in[29]~95 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[29]~96 (
	.dataa(\wb_alu_out[29]~q ),
	.datab(\csr_io_in[0]~2_combout ),
	.datac(\csr_io_in[29]~95_combout ),
	.datad(\wb_csr_data[29]~q ),
	.cin(gnd),
	.combout(\csr_io_in[29]~96_combout ),
	.cout());
defparam \csr_io_in[29]~96 .lut_mask = 16'hF838;
defparam \csr_io_in[29]~96 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[29]~97 (
	.dataa(\mem_csr_data[29]~q ),
	.datab(\csr_io_in[29]~96_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[29]~97_combout ),
	.cout());
defparam \csr_io_in[29]~97 .lut_mask = 16'h00AC;
defparam \csr_io_in[29]~97 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[30]~98 (
	.dataa(\csr_io_in[0]~1_combout ),
	.datab(\wb_alu_out[30]~q ),
	.datac(\csr_io_in[0]~2_combout ),
	.datad(\ex_reg_rs1_bypass[30]~29_combout ),
	.cin(gnd),
	.combout(\csr_io_in[30]~98_combout ),
	.cout());
defparam \csr_io_in[30]~98 .lut_mask = 16'hE5E0;
defparam \csr_io_in[30]~98 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[30]~99 (
	.dataa(\mem_alu_out[30]~q ),
	.datab(\csr_io_in[0]~1_combout ),
	.datac(\csr_io_in[30]~98_combout ),
	.datad(\wb_csr_data[30]~q ),
	.cin(gnd),
	.combout(\csr_io_in[30]~99_combout ),
	.cout());
defparam \csr_io_in[30]~99 .lut_mask = 16'hF838;
defparam \csr_io_in[30]~99 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[30]~100 (
	.dataa(\mem_csr_data[30]~q ),
	.datab(\csr_io_in[30]~99_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[30]~100_combout ),
	.cout());
defparam \csr_io_in[30]~100 .lut_mask = 16'h00AC;
defparam \csr_io_in[30]~100 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[31]~101 (
	.dataa(\wb_csr_data[31]~q ),
	.datab(\wb_alu_out[31]~q ),
	.datac(gnd),
	.datad(\wb_ctrl_csr_cmd.000~q ),
	.cin(gnd),
	.combout(\csr_io_in[31]~101_combout ),
	.cout());
defparam \csr_io_in[31]~101 .lut_mask = 16'hAACC;
defparam \csr_io_in[31]~101 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[31]~102 (
	.dataa(\csr_io_in[31]~101_combout ),
	.datab(\ex_reg_rs1_bypass[31]~33_combout ),
	.datac(\Equal61~2_combout ),
	.datad(\Equal60~5_combout ),
	.cin(gnd),
	.combout(\csr_io_in[31]~102_combout ),
	.cout());
defparam \csr_io_in[31]~102 .lut_mask = 16'h00AC;
defparam \csr_io_in[31]~102 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[31]~103 (
	.dataa(\mem_csr_data[31]~q ),
	.datab(\mem_alu_out[31]~q ),
	.datac(gnd),
	.datad(\mem_ctrl_csr_cmd.000~q ),
	.cin(gnd),
	.combout(\csr_io_in[31]~103_combout ),
	.cout());
defparam \csr_io_in[31]~103 .lut_mask = 16'hAACC;
defparam \csr_io_in[31]~103 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[31]~104 (
	.dataa(\csr_io_in[31]~102_combout ),
	.datab(\Equal60~5_combout ),
	.datac(\csr_io_in[31]~103_combout ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\csr_io_in[31]~104_combout ),
	.cout());
defparam \csr_io_in[31]~104 .lut_mask = 16'h00EA;
defparam \csr_io_in[31]~104 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_inst~13 (
	.dataa(\id_inst[0]~q ),
	.datab(gnd),
	.datac(\_T_1778~combout ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\ex_inst~13_combout ),
	.cout());
defparam \ex_inst~13 .lut_mask = 16'hAFFF;
defparam \ex_inst~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_inst~14 (
	.dataa(\id_inst[1]~q ),
	.datab(gnd),
	.datac(\_T_1778~combout ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\ex_inst~14_combout ),
	.cout());
defparam \ex_inst~14 .lut_mask = 16'hAFFF;
defparam \ex_inst~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_inst~15 (
	.dataa(\id_inst[4]~q ),
	.datab(gnd),
	.datac(\_T_1778~combout ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\ex_inst~15_combout ),
	.cout());
defparam \ex_inst~15 .lut_mask = 16'hAFFF;
defparam \ex_inst~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_inst~16 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~16_combout ),
	.cout());
defparam \ex_inst~16 .lut_mask = 16'h8080;
defparam \ex_inst~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_inst~17 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~17_combout ),
	.cout());
defparam \ex_inst~17 .lut_mask = 16'h8080;
defparam \ex_inst~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_inst~18 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~18_combout ),
	.cout());
defparam \ex_inst~18 .lut_mask = 16'h8080;
defparam \ex_inst~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_inst~19 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[6]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~19_combout ),
	.cout());
defparam \ex_inst~19 .lut_mask = 16'h8080;
defparam \ex_inst~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_legal~3 (
	.dataa(\Equal53~0_combout ),
	.datab(\Equal18~0_combout ),
	.datac(\id_inst[14]~q ),
	.datad(\id_inst[4]~q ),
	.cin(gnd),
	.combout(\ex_ctrl_legal~3_combout ),
	.cout());
defparam \ex_ctrl_legal~3 .lut_mask = 16'h0008;
defparam \ex_ctrl_legal~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_GEN_33~2 (
	.dataa(\id_inst[12]~q ),
	.datab(\Equal11~0_combout ),
	.datac(\id_ctrl_br_type[2]~5_combout ),
	.datad(\_T_1778~combout ),
	.cin(gnd),
	.combout(\_GEN_33~2_combout ),
	.cout());
defparam \_GEN_33~2 .lut_mask = 16'hF400;
defparam \_GEN_33~2 .sum_lutc_input = "datac";

dffeas \id_npc[0] (
	.clk(clk_clk),
	.d(\id_npc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_npc_0),
	.prn(vcc));
defparam \id_npc[0] .is_wysiwyg = "true";
defparam \id_npc[0] .power_up = "low";

dffeas \id_npc[1] (
	.clk(clk_clk),
	.d(\id_npc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_npc_1),
	.prn(vcc));
defparam \id_npc[1] .is_wysiwyg = "true";
defparam \id_npc[1] .power_up = "low";

dffeas \id_pc[2] (
	.clk(clk_clk),
	.d(\id_pc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_2),
	.prn(vcc));
defparam \id_pc[2] .is_wysiwyg = "true";
defparam \id_pc[2] .power_up = "low";

dffeas \id_pc[3] (
	.clk(clk_clk),
	.d(\id_pc~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_3),
	.prn(vcc));
defparam \id_pc[3] .is_wysiwyg = "true";
defparam \id_pc[3] .power_up = "low";

dffeas \id_pc[4] (
	.clk(clk_clk),
	.d(\id_pc~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_4),
	.prn(vcc));
defparam \id_pc[4] .is_wysiwyg = "true";
defparam \id_pc[4] .power_up = "low";

dffeas \id_pc[5] (
	.clk(clk_clk),
	.d(\id_pc~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_5),
	.prn(vcc));
defparam \id_pc[5] .is_wysiwyg = "true";
defparam \id_pc[5] .power_up = "low";

dffeas \id_pc[6] (
	.clk(clk_clk),
	.d(\id_pc~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_6),
	.prn(vcc));
defparam \id_pc[6] .is_wysiwyg = "true";
defparam \id_pc[6] .power_up = "low";

dffeas \id_pc[7] (
	.clk(clk_clk),
	.d(\id_pc~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_7),
	.prn(vcc));
defparam \id_pc[7] .is_wysiwyg = "true";
defparam \id_pc[7] .power_up = "low";

dffeas \id_pc[8] (
	.clk(clk_clk),
	.d(\id_pc~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_8),
	.prn(vcc));
defparam \id_pc[8] .is_wysiwyg = "true";
defparam \id_pc[8] .power_up = "low";

dffeas \id_pc[9] (
	.clk(clk_clk),
	.d(\id_pc~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_9),
	.prn(vcc));
defparam \id_pc[9] .is_wysiwyg = "true";
defparam \id_pc[9] .power_up = "low";

dffeas \id_pc[10] (
	.clk(clk_clk),
	.d(\id_pc~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_10),
	.prn(vcc));
defparam \id_pc[10] .is_wysiwyg = "true";
defparam \id_pc[10] .power_up = "low";

dffeas \id_pc[11] (
	.clk(clk_clk),
	.d(\id_pc~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_11),
	.prn(vcc));
defparam \id_pc[11] .is_wysiwyg = "true";
defparam \id_pc[11] .power_up = "low";

dffeas \id_pc[12] (
	.clk(clk_clk),
	.d(\id_pc~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_12),
	.prn(vcc));
defparam \id_pc[12] .is_wysiwyg = "true";
defparam \id_pc[12] .power_up = "low";

dffeas \id_pc[13] (
	.clk(clk_clk),
	.d(\id_pc~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_13),
	.prn(vcc));
defparam \id_pc[13] .is_wysiwyg = "true";
defparam \id_pc[13] .power_up = "low";

dffeas \id_pc[14] (
	.clk(clk_clk),
	.d(\id_pc~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_14),
	.prn(vcc));
defparam \id_pc[14] .is_wysiwyg = "true";
defparam \id_pc[14] .power_up = "low";

dffeas \id_pc[15] (
	.clk(clk_clk),
	.d(\id_pc~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_15),
	.prn(vcc));
defparam \id_pc[15] .is_wysiwyg = "true";
defparam \id_pc[15] .power_up = "low";

dffeas \id_pc[16] (
	.clk(clk_clk),
	.d(\id_pc~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_16),
	.prn(vcc));
defparam \id_pc[16] .is_wysiwyg = "true";
defparam \id_pc[16] .power_up = "low";

dffeas \id_pc[17] (
	.clk(clk_clk),
	.d(\id_pc~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_17),
	.prn(vcc));
defparam \id_pc[17] .is_wysiwyg = "true";
defparam \id_pc[17] .power_up = "low";

dffeas \id_pc[18] (
	.clk(clk_clk),
	.d(\id_pc~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_18),
	.prn(vcc));
defparam \id_pc[18] .is_wysiwyg = "true";
defparam \id_pc[18] .power_up = "low";

dffeas \id_pc[19] (
	.clk(clk_clk),
	.d(\id_pc~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_19),
	.prn(vcc));
defparam \id_pc[19] .is_wysiwyg = "true";
defparam \id_pc[19] .power_up = "low";

dffeas \id_pc[20] (
	.clk(clk_clk),
	.d(\id_pc~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_20),
	.prn(vcc));
defparam \id_pc[20] .is_wysiwyg = "true";
defparam \id_pc[20] .power_up = "low";

dffeas \id_pc[21] (
	.clk(clk_clk),
	.d(\id_pc~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_21),
	.prn(vcc));
defparam \id_pc[21] .is_wysiwyg = "true";
defparam \id_pc[21] .power_up = "low";

dffeas \id_pc[22] (
	.clk(clk_clk),
	.d(\id_pc~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_22),
	.prn(vcc));
defparam \id_pc[22] .is_wysiwyg = "true";
defparam \id_pc[22] .power_up = "low";

dffeas \id_pc[23] (
	.clk(clk_clk),
	.d(\id_pc~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_23),
	.prn(vcc));
defparam \id_pc[23] .is_wysiwyg = "true";
defparam \id_pc[23] .power_up = "low";

dffeas \id_pc[24] (
	.clk(clk_clk),
	.d(\id_pc~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_24),
	.prn(vcc));
defparam \id_pc[24] .is_wysiwyg = "true";
defparam \id_pc[24] .power_up = "low";

dffeas \id_pc[25] (
	.clk(clk_clk),
	.d(\id_pc~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_25),
	.prn(vcc));
defparam \id_pc[25] .is_wysiwyg = "true";
defparam \id_pc[25] .power_up = "low";

dffeas \id_pc[26] (
	.clk(clk_clk),
	.d(\id_pc~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_26),
	.prn(vcc));
defparam \id_pc[26] .is_wysiwyg = "true";
defparam \id_pc[26] .power_up = "low";

dffeas \id_pc[27] (
	.clk(clk_clk),
	.d(\id_pc~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_27),
	.prn(vcc));
defparam \id_pc[27] .is_wysiwyg = "true";
defparam \id_pc[27] .power_up = "low";

dffeas \id_pc[28] (
	.clk(clk_clk),
	.d(\id_pc~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_28),
	.prn(vcc));
defparam \id_pc[28] .is_wysiwyg = "true";
defparam \id_pc[28] .power_up = "low";

dffeas \id_pc[29] (
	.clk(clk_clk),
	.d(\id_pc~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_29),
	.prn(vcc));
defparam \id_pc[29] .is_wysiwyg = "true";
defparam \id_pc[29] .power_up = "low";

dffeas \id_pc[30] (
	.clk(clk_clk),
	.d(\id_pc~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_30),
	.prn(vcc));
defparam \id_pc[30] .is_wysiwyg = "true";
defparam \id_pc[30] .power_up = "low";

dffeas \id_pc[31] (
	.clk(clk_clk),
	.d(\id_pc~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(id_pc_31),
	.prn(vcc));
defparam \id_pc[31] .is_wysiwyg = "true";
defparam \id_pc[31] .power_up = "low";

dffeas \mem_alu_out[1] (
	.clk(clk_clk),
	.d(\mem_alu_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_alu_out_1),
	.prn(vcc));
defparam \mem_alu_out[1] .is_wysiwyg = "true";
defparam \mem_alu_out[1] .power_up = "low";

dffeas \mem_alu_out[0] (
	.clk(clk_clk),
	.d(\mem_alu_out~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_alu_out_0),
	.prn(vcc));
defparam \mem_alu_out[0] .is_wysiwyg = "true";
defparam \mem_alu_out[0] .power_up = "low";

dffeas \mem_ctrl_mem_wr.10 (
	.clk(clk_clk),
	.d(\mem_ctrl_mem_wr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_ctrl_mem_wr10),
	.prn(vcc));
defparam \mem_ctrl_mem_wr.10 .is_wysiwyg = "true";
defparam \mem_ctrl_mem_wr.10 .power_up = "low";

dffeas \mem_rs_1[0] (
	.clk(clk_clk),
	.d(\mem_rs_1~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_0),
	.prn(vcc));
defparam \mem_rs_1[0] .is_wysiwyg = "true";
defparam \mem_rs_1[0] .power_up = "low";

cyclone10lp_lcell_comb \Equal68~0 (
	.dataa(\mem_ctrl_mask_type[0]~q ),
	.datab(gnd),
	.datac(\mem_ctrl_mask_type[2]~q ),
	.datad(\mem_ctrl_mask_type[1]~q ),
	.cin(gnd),
	.combout(Equal68),
	.cout());
defparam \Equal68~0 .lut_mask = 16'h000A;
defparam \Equal68~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal73~0 (
	.dataa(\mem_ctrl_mask_type[1]~q ),
	.datab(gnd),
	.datac(\mem_ctrl_mask_type[2]~q ),
	.datad(\mem_ctrl_mask_type[0]~q ),
	.cin(gnd),
	.combout(Equal73),
	.cout());
defparam \Equal73~0 .lut_mask = 16'h000A;
defparam \Equal73~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[0]~16 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(mem_rs_1_0),
	.datac(_GEN_73_0),
	.datad(gnd),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_0),
	.cout());
defparam \io_w_dmem_dat_data[0]~16 .lut_mask = 16'h8080;
defparam \io_w_dmem_dat_data[0]~16 .sum_lutc_input = "datac";

dffeas \mem_alu_out[2] (
	.clk(clk_clk),
	.d(\mem_alu_out~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_alu_out_2),
	.prn(vcc));
defparam \mem_alu_out[2] .is_wysiwyg = "true";
defparam \mem_alu_out[2] .power_up = "low";

dffeas \mem_alu_out[3] (
	.clk(clk_clk),
	.d(\mem_alu_out~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_alu_out_3),
	.prn(vcc));
defparam \mem_alu_out[3] .is_wysiwyg = "true";
defparam \mem_alu_out[3] .power_up = "low";

dffeas \mem_rs_1[1] (
	.clk(clk_clk),
	.d(\mem_rs_1~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_1),
	.prn(vcc));
defparam \mem_rs_1[1] .is_wysiwyg = "true";
defparam \mem_rs_1[1] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[1]~17 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(_GEN_73_0),
	.datac(mem_rs_1_1),
	.datad(gnd),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_1),
	.cout());
defparam \io_w_dmem_dat_data[1]~17 .lut_mask = 16'h8080;
defparam \io_w_dmem_dat_data[1]~17 .sum_lutc_input = "datac";

dffeas \mem_rs_1[2] (
	.clk(clk_clk),
	.d(\mem_rs_1~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_2),
	.prn(vcc));
defparam \mem_rs_1[2] .is_wysiwyg = "true";
defparam \mem_rs_1[2] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[2]~18 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(_GEN_73_0),
	.datac(mem_rs_1_2),
	.datad(gnd),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_2),
	.cout());
defparam \io_w_dmem_dat_data[2]~18 .lut_mask = 16'h8080;
defparam \io_w_dmem_dat_data[2]~18 .sum_lutc_input = "datac";

dffeas \mem_rs_1[3] (
	.clk(clk_clk),
	.d(\mem_rs_1~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_3),
	.prn(vcc));
defparam \mem_rs_1[3] .is_wysiwyg = "true";
defparam \mem_rs_1[3] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[3]~19 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(_GEN_73_0),
	.datac(mem_rs_1_3),
	.datad(gnd),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_3),
	.cout());
defparam \io_w_dmem_dat_data[3]~19 .lut_mask = 16'h8080;
defparam \io_w_dmem_dat_data[3]~19 .sum_lutc_input = "datac";

dffeas \mem_rs_1[4] (
	.clk(clk_clk),
	.d(\mem_rs_1~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_4),
	.prn(vcc));
defparam \mem_rs_1[4] .is_wysiwyg = "true";
defparam \mem_rs_1[4] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[4]~20 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(_GEN_73_0),
	.datac(mem_rs_1_4),
	.datad(gnd),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_4),
	.cout());
defparam \io_w_dmem_dat_data[4]~20 .lut_mask = 16'h8080;
defparam \io_w_dmem_dat_data[4]~20 .sum_lutc_input = "datac";

dffeas \mem_rs_1[5] (
	.clk(clk_clk),
	.d(\mem_rs_1~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_5),
	.prn(vcc));
defparam \mem_rs_1[5] .is_wysiwyg = "true";
defparam \mem_rs_1[5] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[5]~21 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(_GEN_73_0),
	.datac(mem_rs_1_5),
	.datad(gnd),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_5),
	.cout());
defparam \io_w_dmem_dat_data[5]~21 .lut_mask = 16'h8080;
defparam \io_w_dmem_dat_data[5]~21 .sum_lutc_input = "datac";

dffeas \mem_rs_1[6] (
	.clk(clk_clk),
	.d(\mem_rs_1~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_6),
	.prn(vcc));
defparam \mem_rs_1[6] .is_wysiwyg = "true";
defparam \mem_rs_1[6] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[6]~22 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(_GEN_73_0),
	.datac(mem_rs_1_6),
	.datad(gnd),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_6),
	.cout());
defparam \io_w_dmem_dat_data[6]~22 .lut_mask = 16'h8080;
defparam \io_w_dmem_dat_data[6]~22 .sum_lutc_input = "datac";

dffeas \mem_rs_1[7] (
	.clk(clk_clk),
	.d(\mem_rs_1~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_7),
	.prn(vcc));
defparam \mem_rs_1[7] .is_wysiwyg = "true";
defparam \mem_rs_1[7] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[7]~23 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(_GEN_73_0),
	.datac(mem_rs_1_7),
	.datad(gnd),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_7),
	.cout());
defparam \io_w_dmem_dat_data[7]~23 .lut_mask = 16'h8080;
defparam \io_w_dmem_dat_data[7]~23 .sum_lutc_input = "datac";

dffeas \mem_rs_1[8] (
	.clk(clk_clk),
	.d(\mem_rs_1~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_8),
	.prn(vcc));
defparam \mem_rs_1[8] .is_wysiwyg = "true";
defparam \mem_rs_1[8] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[8]~24 (
	.dataa(mem_rs_1_8),
	.datab(mem_rs_1_0),
	.datac(_GEN_73_0),
	.datad(data_out_12),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_8),
	.cout());
defparam \io_w_dmem_dat_data[8]~24 .lut_mask = 16'h00AC;
defparam \io_w_dmem_dat_data[8]~24 .sum_lutc_input = "datac";

dffeas \mem_rs_1[9] (
	.clk(clk_clk),
	.d(\mem_rs_1~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_9),
	.prn(vcc));
defparam \mem_rs_1[9] .is_wysiwyg = "true";
defparam \mem_rs_1[9] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[9]~25 (
	.dataa(mem_rs_1_9),
	.datab(mem_rs_1_1),
	.datac(_GEN_73_0),
	.datad(data_out_12),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_9),
	.cout());
defparam \io_w_dmem_dat_data[9]~25 .lut_mask = 16'h00AC;
defparam \io_w_dmem_dat_data[9]~25 .sum_lutc_input = "datac";

dffeas \mem_rs_1[10] (
	.clk(clk_clk),
	.d(\mem_rs_1~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_10),
	.prn(vcc));
defparam \mem_rs_1[10] .is_wysiwyg = "true";
defparam \mem_rs_1[10] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[10]~26 (
	.dataa(mem_rs_1_10),
	.datab(mem_rs_1_2),
	.datac(_GEN_73_0),
	.datad(data_out_12),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_10),
	.cout());
defparam \io_w_dmem_dat_data[10]~26 .lut_mask = 16'h00AC;
defparam \io_w_dmem_dat_data[10]~26 .sum_lutc_input = "datac";

dffeas \mem_rs_1[11] (
	.clk(clk_clk),
	.d(\mem_rs_1~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_11),
	.prn(vcc));
defparam \mem_rs_1[11] .is_wysiwyg = "true";
defparam \mem_rs_1[11] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[11]~27 (
	.dataa(mem_rs_1_11),
	.datab(mem_rs_1_3),
	.datac(_GEN_73_0),
	.datad(data_out_12),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_11),
	.cout());
defparam \io_w_dmem_dat_data[11]~27 .lut_mask = 16'h00AC;
defparam \io_w_dmem_dat_data[11]~27 .sum_lutc_input = "datac";

dffeas \mem_rs_1[12] (
	.clk(clk_clk),
	.d(\mem_rs_1~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_12),
	.prn(vcc));
defparam \mem_rs_1[12] .is_wysiwyg = "true";
defparam \mem_rs_1[12] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[12]~28 (
	.dataa(mem_rs_1_12),
	.datab(mem_rs_1_4),
	.datac(_GEN_73_0),
	.datad(data_out_12),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_12),
	.cout());
defparam \io_w_dmem_dat_data[12]~28 .lut_mask = 16'h00AC;
defparam \io_w_dmem_dat_data[12]~28 .sum_lutc_input = "datac";

dffeas \mem_rs_1[13] (
	.clk(clk_clk),
	.d(\mem_rs_1~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_13),
	.prn(vcc));
defparam \mem_rs_1[13] .is_wysiwyg = "true";
defparam \mem_rs_1[13] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[13]~29 (
	.dataa(mem_rs_1_13),
	.datab(mem_rs_1_5),
	.datac(_GEN_73_0),
	.datad(data_out_12),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_13),
	.cout());
defparam \io_w_dmem_dat_data[13]~29 .lut_mask = 16'h00AC;
defparam \io_w_dmem_dat_data[13]~29 .sum_lutc_input = "datac";

dffeas \mem_rs_1[14] (
	.clk(clk_clk),
	.d(\mem_rs_1~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_14),
	.prn(vcc));
defparam \mem_rs_1[14] .is_wysiwyg = "true";
defparam \mem_rs_1[14] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[14]~30 (
	.dataa(mem_rs_1_14),
	.datab(mem_rs_1_6),
	.datac(_GEN_73_0),
	.datad(data_out_12),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_14),
	.cout());
defparam \io_w_dmem_dat_data[14]~30 .lut_mask = 16'h00AC;
defparam \io_w_dmem_dat_data[14]~30 .sum_lutc_input = "datac";

dffeas \mem_rs_1[15] (
	.clk(clk_clk),
	.d(\mem_rs_1~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_15),
	.prn(vcc));
defparam \mem_rs_1[15] .is_wysiwyg = "true";
defparam \mem_rs_1[15] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[15]~31 (
	.dataa(mem_rs_1_15),
	.datab(mem_rs_1_7),
	.datac(_GEN_73_0),
	.datad(data_out_12),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_15),
	.cout());
defparam \io_w_dmem_dat_data[15]~31 .lut_mask = 16'h00AC;
defparam \io_w_dmem_dat_data[15]~31 .sum_lutc_input = "datac";

dffeas \mem_rs_1[16] (
	.clk(clk_clk),
	.d(\mem_rs_1~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_16),
	.prn(vcc));
defparam \mem_rs_1[16] .is_wysiwyg = "true";
defparam \mem_rs_1[16] .power_up = "low";

dffeas \mem_rs_1[17] (
	.clk(clk_clk),
	.d(\mem_rs_1~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_17),
	.prn(vcc));
defparam \mem_rs_1[17] .is_wysiwyg = "true";
defparam \mem_rs_1[17] .power_up = "low";

dffeas \mem_rs_1[18] (
	.clk(clk_clk),
	.d(\mem_rs_1~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_18),
	.prn(vcc));
defparam \mem_rs_1[18] .is_wysiwyg = "true";
defparam \mem_rs_1[18] .power_up = "low";

dffeas \mem_rs_1[19] (
	.clk(clk_clk),
	.d(\mem_rs_1~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_19),
	.prn(vcc));
defparam \mem_rs_1[19] .is_wysiwyg = "true";
defparam \mem_rs_1[19] .power_up = "low";

dffeas \mem_rs_1[20] (
	.clk(clk_clk),
	.d(\mem_rs_1~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_20),
	.prn(vcc));
defparam \mem_rs_1[20] .is_wysiwyg = "true";
defparam \mem_rs_1[20] .power_up = "low";

dffeas \mem_rs_1[21] (
	.clk(clk_clk),
	.d(\mem_rs_1~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_21),
	.prn(vcc));
defparam \mem_rs_1[21] .is_wysiwyg = "true";
defparam \mem_rs_1[21] .power_up = "low";

dffeas \mem_rs_1[22] (
	.clk(clk_clk),
	.d(\mem_rs_1~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_22),
	.prn(vcc));
defparam \mem_rs_1[22] .is_wysiwyg = "true";
defparam \mem_rs_1[22] .power_up = "low";

dffeas \mem_rs_1[23] (
	.clk(clk_clk),
	.d(\mem_rs_1~65_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rs_1_23),
	.prn(vcc));
defparam \mem_rs_1[23] .is_wysiwyg = "true";
defparam \mem_rs_1[23] .power_up = "low";

dffeas \mem_ctrl_mem_wr.00 (
	.clk(clk_clk),
	.d(\mem_ctrl_mem_wr~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_ctrl_mem_wr00),
	.prn(vcc));
defparam \mem_ctrl_mem_wr.00 .is_wysiwyg = "true";
defparam \mem_ctrl_mem_wr.00 .power_up = "low";

dffeas w_req(
	.clk(clk_clk),
	.d(\w_req~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(w_req1),
	.prn(vcc));
defparam w_req.is_wysiwyg = "true";
defparam w_req.power_up = "low";

dffeas \mem_ctrl_mem_wr.01 (
	.clk(clk_clk),
	.d(\mem_ctrl_mem_wr~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_ctrl_mem_wr01),
	.prn(vcc));
defparam \mem_ctrl_mem_wr.01 .is_wysiwyg = "true";
defparam \mem_ctrl_mem_wr.01 .power_up = "low";

cyclone10lp_lcell_comb \io_imem_add_addr[2]~0 (
	.dataa(\pc_cntr[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(w_req1),
	.cin(gnd),
	.combout(io_imem_add_addr_2),
	.cout());
defparam \io_imem_add_addr[2]~0 .lut_mask = 16'h00AA;
defparam \io_imem_add_addr[2]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_imem_add_addr[3]~1 (
	.dataa(\pc_cntr[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(w_req1),
	.cin(gnd),
	.combout(io_imem_add_addr_3),
	.cout());
defparam \io_imem_add_addr[3]~1 .lut_mask = 16'h00AA;
defparam \io_imem_add_addr[3]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_imem_add_addr[4]~2 (
	.dataa(\pc_cntr[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(w_req1),
	.cin(gnd),
	.combout(io_imem_add_addr_4),
	.cout());
defparam \io_imem_add_addr[4]~2 .lut_mask = 16'h00AA;
defparam \io_imem_add_addr[4]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_imem_add_addr[5]~3 (
	.dataa(\pc_cntr[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(w_req1),
	.cin(gnd),
	.combout(io_imem_add_addr_5),
	.cout());
defparam \io_imem_add_addr[5]~3 .lut_mask = 16'h00AA;
defparam \io_imem_add_addr[5]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_imem_add_addr[6]~4 (
	.dataa(\pc_cntr[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(w_req1),
	.cin(gnd),
	.combout(io_imem_add_addr_6),
	.cout());
defparam \io_imem_add_addr[6]~4 .lut_mask = 16'h00AA;
defparam \io_imem_add_addr[6]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_imem_add_addr[7]~5 (
	.dataa(\pc_cntr[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(w_req1),
	.cin(gnd),
	.combout(io_imem_add_addr_7),
	.cout());
defparam \io_imem_add_addr[7]~5 .lut_mask = 16'h00AA;
defparam \io_imem_add_addr[7]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_imem_add_addr[8]~6 (
	.dataa(\pc_cntr[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(w_req1),
	.cin(gnd),
	.combout(io_imem_add_addr_8),
	.cout());
defparam \io_imem_add_addr[8]~6 .lut_mask = 16'h00AA;
defparam \io_imem_add_addr[8]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_imem_add_addr[9]~7 (
	.dataa(\pc_cntr[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(w_req1),
	.cin(gnd),
	.combout(io_imem_add_addr_9),
	.cout());
defparam \io_imem_add_addr[9]~7 .lut_mask = 16'h00AA;
defparam \io_imem_add_addr[9]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_imem_add_addr[10]~8 (
	.dataa(\pc_cntr[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(w_req1),
	.cin(gnd),
	.combout(io_imem_add_addr_10),
	.cout());
defparam \io_imem_add_addr[10]~8 .lut_mask = 16'h00AA;
defparam \io_imem_add_addr[10]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_imem_add_addr[11]~9 (
	.dataa(\pc_cntr[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(w_req1),
	.cin(gnd),
	.combout(io_imem_add_addr_11),
	.cout());
defparam \io_imem_add_addr[11]~9 .lut_mask = 16'h00AA;
defparam \io_imem_add_addr[11]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_imem_add_addr[12]~10 (
	.dataa(\pc_cntr[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(w_req1),
	.cin(gnd),
	.combout(io_imem_add_addr_12),
	.cout());
defparam \io_imem_add_addr[12]~10 .lut_mask = 16'h00AA;
defparam \io_imem_add_addr[12]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_imem_add_addr[13]~11 (
	.dataa(\pc_cntr[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(w_req1),
	.cin(gnd),
	.combout(io_imem_add_addr_13),
	.cout());
defparam \io_imem_add_addr[13]~11 .lut_mask = 16'h00AA;
defparam \io_imem_add_addr[13]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_imem_add_addr[14]~12 (
	.dataa(\pc_cntr[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(w_req1),
	.cin(gnd),
	.combout(io_imem_add_addr_14),
	.cout());
defparam \io_imem_add_addr[14]~12 .lut_mask = 16'h00AA;
defparam \io_imem_add_addr[14]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_GEN_73[0]~2 (
	.dataa(mem_alu_out_0),
	.datab(mem_alu_out_1),
	.datac(Equal68),
	.datad(Equal73),
	.cin(gnd),
	.combout(_GEN_73_0),
	.cout());
defparam \_GEN_73[0]~2 .lut_mask = 16'h111F;
defparam \_GEN_73[0]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[24]~48 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(mem_alu_out_0),
	.datac(Equal73),
	.datad(\io_w_dmem_dat_data[24]~33_combout ),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_24),
	.cout());
defparam \io_w_dmem_dat_data[24]~48 .lut_mask = 16'h2A00;
defparam \io_w_dmem_dat_data[24]~48 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[25]~49 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(mem_alu_out_0),
	.datac(Equal73),
	.datad(\io_w_dmem_dat_data[25]~35_combout ),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_25),
	.cout());
defparam \io_w_dmem_dat_data[25]~49 .lut_mask = 16'h2A00;
defparam \io_w_dmem_dat_data[25]~49 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[26]~50 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(mem_alu_out_0),
	.datac(Equal73),
	.datad(\io_w_dmem_dat_data[26]~37_combout ),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_26),
	.cout());
defparam \io_w_dmem_dat_data[26]~50 .lut_mask = 16'h2A00;
defparam \io_w_dmem_dat_data[26]~50 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[27]~51 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(mem_alu_out_0),
	.datac(Equal73),
	.datad(\io_w_dmem_dat_data[27]~39_combout ),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_27),
	.cout());
defparam \io_w_dmem_dat_data[27]~51 .lut_mask = 16'h2A00;
defparam \io_w_dmem_dat_data[27]~51 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[28]~52 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(mem_alu_out_0),
	.datac(Equal73),
	.datad(\io_w_dmem_dat_data[28]~41_combout ),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_28),
	.cout());
defparam \io_w_dmem_dat_data[28]~52 .lut_mask = 16'h2A00;
defparam \io_w_dmem_dat_data[28]~52 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[29]~53 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(mem_alu_out_0),
	.datac(Equal73),
	.datad(\io_w_dmem_dat_data[29]~43_combout ),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_29),
	.cout());
defparam \io_w_dmem_dat_data[29]~53 .lut_mask = 16'h2A00;
defparam \io_w_dmem_dat_data[29]~53 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[30]~54 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(mem_alu_out_0),
	.datac(Equal73),
	.datad(\io_w_dmem_dat_data[30]~45_combout ),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_30),
	.cout());
defparam \io_w_dmem_dat_data[30]~54 .lut_mask = 16'h2A00;
defparam \io_w_dmem_dat_data[30]~54 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[31]~55 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(mem_alu_out_0),
	.datac(Equal73),
	.datad(\io_w_dmem_dat_data[31]~47_combout ),
	.cin(gnd),
	.combout(io_w_dmem_dat_data_31),
	.cout());
defparam \io_w_dmem_dat_data[31]~55 .lut_mask = 16'h2A00;
defparam \io_w_dmem_dat_data[31]~55 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb _T_1778(
	.dataa(\inst_kill~0_combout ),
	.datab(\csr|io_expt~0_combout ),
	.datac(\csr|mcause[0]~6_combout ),
	.datad(\csr|isEcall~0_combout ),
	.cin(gnd),
	.combout(\_T_1778~combout ),
	.cout());
defparam _T_1778.lut_mask = 16'h0080;
defparam _T_1778.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~21 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_14),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~21_combout ),
	.cout());
defparam \id_inst~21 .lut_mask = 16'h8080;
defparam \id_inst~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~0 (
	.dataa(\inst_kill~0_combout ),
	.datab(\csr|io_expt~0_combout ),
	.datac(\csr|isEcall~0_combout ),
	.datad(\csr|mcause[0]~6_combout ),
	.cin(gnd),
	.combout(\id_inst~0_combout ),
	.cout());
defparam \id_inst~0 .lut_mask = 16'h0008;
defparam \id_inst~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_pc[7]~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\id_inst~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc[7]~0_combout ),
	.cout());
defparam \id_pc[7]~0 .lut_mask = 16'h7777;
defparam \id_pc[7]~0 .sum_lutc_input = "datac";

dffeas \id_inst[14] (
	.clk(clk_clk),
	.d(\id_inst~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[14]~q ),
	.prn(vcc));
defparam \id_inst[14] .is_wysiwyg = "true";
defparam \id_inst[14] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~33 (
	.dataa(q_a_0),
	.datab(gnd),
	.datac(\_T_1778~combout ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\id_inst~33_combout ),
	.cout());
defparam \id_inst~33 .lut_mask = 16'hAFFF;
defparam \id_inst~33 .sum_lutc_input = "datac";

dffeas \id_inst[0] (
	.clk(clk_clk),
	.d(\id_inst~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[0]~q ),
	.prn(vcc));
defparam \id_inst[0] .is_wysiwyg = "true";
defparam \id_inst[0] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~34 (
	.dataa(q_a_1),
	.datab(gnd),
	.datac(\_T_1778~combout ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\id_inst~34_combout ),
	.cout());
defparam \id_inst~34 .lut_mask = 16'hAFFF;
defparam \id_inst~34 .sum_lutc_input = "datac";

dffeas \id_inst[1] (
	.clk(clk_clk),
	.d(\id_inst~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[1]~q ),
	.prn(vcc));
defparam \id_inst[1] .is_wysiwyg = "true";
defparam \id_inst[1] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~35 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_3),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~35_combout ),
	.cout());
defparam \id_inst~35 .lut_mask = 16'h8080;
defparam \id_inst~35 .sum_lutc_input = "datac";

dffeas \id_inst[3] (
	.clk(clk_clk),
	.d(\id_inst~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[3]~q ),
	.prn(vcc));
defparam \id_inst[3] .is_wysiwyg = "true";
defparam \id_inst[3] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~36 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~36_combout ),
	.cout());
defparam \id_inst~36 .lut_mask = 16'h8080;
defparam \id_inst~36 .sum_lutc_input = "datac";

dffeas \id_inst[2] (
	.clk(clk_clk),
	.d(\id_inst~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[2]~q ),
	.prn(vcc));
defparam \id_inst[2] .is_wysiwyg = "true";
defparam \id_inst[2] .power_up = "low";

cyclone10lp_lcell_comb \ex_ctrl_mem_wr~7 (
	.dataa(\id_inst[0]~q ),
	.datab(\id_inst[1]~q ),
	.datac(\id_inst[3]~q ),
	.datad(\id_inst[2]~q ),
	.cin(gnd),
	.combout(\ex_ctrl_mem_wr~7_combout ),
	.cout());
defparam \ex_ctrl_mem_wr~7 .lut_mask = 16'h0008;
defparam \ex_ctrl_mem_wr~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~23 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_5),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~23_combout ),
	.cout());
defparam \id_inst~23 .lut_mask = 16'h8080;
defparam \id_inst~23 .sum_lutc_input = "datac";

dffeas \id_inst[5] (
	.clk(clk_clk),
	.d(\id_inst~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[5]~q ),
	.prn(vcc));
defparam \id_inst[5] .is_wysiwyg = "true";
defparam \id_inst[5] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~24 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_6),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~24_combout ),
	.cout());
defparam \id_inst~24 .lut_mask = 16'h8080;
defparam \id_inst~24 .sum_lutc_input = "datac";

dffeas \id_inst[6] (
	.clk(clk_clk),
	.d(\id_inst~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[6]~q ),
	.prn(vcc));
defparam \id_inst[6] .is_wysiwyg = "true";
defparam \id_inst[6] .power_up = "low";

cyclone10lp_lcell_comb \Equal7~0 (
	.dataa(\id_inst[5]~q ),
	.datab(\id_inst[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal7~0_combout ),
	.cout());
defparam \Equal7~0 .lut_mask = 16'h8888;
defparam \Equal7~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~37 (
	.dataa(q_a_4),
	.datab(gnd),
	.datac(\_T_1778~combout ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\id_inst~37_combout ),
	.cout());
defparam \id_inst~37 .lut_mask = 16'hAFFF;
defparam \id_inst~37 .sum_lutc_input = "datac";

dffeas \id_inst[4] (
	.clk(clk_clk),
	.d(\id_inst~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[4]~q ),
	.prn(vcc));
defparam \id_inst[4] .is_wysiwyg = "true";
defparam \id_inst[4] .power_up = "low";

cyclone10lp_lcell_comb \Equal11~0 (
	.dataa(\id_inst[14]~q ),
	.datab(\ex_ctrl_mem_wr~7_combout ),
	.datac(\Equal7~0_combout ),
	.datad(\id_inst[4]~q ),
	.cin(gnd),
	.combout(\Equal11~0_combout ),
	.cout());
defparam \Equal11~0 .lut_mask = 16'h0080;
defparam \Equal11~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~28 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_12),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~28_combout ),
	.cout());
defparam \id_inst~28 .lut_mask = 16'h8080;
defparam \id_inst~28 .sum_lutc_input = "datac";

dffeas \id_inst[12] (
	.clk(clk_clk),
	.d(\id_inst~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[12]~q ),
	.prn(vcc));
defparam \id_inst[12] .is_wysiwyg = "true";
defparam \id_inst[12] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~22 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_13),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~22_combout ),
	.cout());
defparam \id_inst~22 .lut_mask = 16'h8080;
defparam \id_inst~22 .sum_lutc_input = "datac";

dffeas \id_inst[13] (
	.clk(clk_clk),
	.d(\id_inst~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[13]~q ),
	.prn(vcc));
defparam \id_inst[13] .is_wysiwyg = "true";
defparam \id_inst[13] .power_up = "low";

cyclone10lp_lcell_comb \Equal14~0 (
	.dataa(\Equal11~0_combout ),
	.datab(\id_inst[12]~q ),
	.datac(\id_inst[13]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal14~0_combout ),
	.cout());
defparam \Equal14~0 .lut_mask = 16'h8080;
defparam \Equal14~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal9~0 (
	.dataa(\ex_ctrl_mem_wr~7_combout ),
	.datab(gnd),
	.datac(\id_inst[14]~q ),
	.datad(\id_inst[13]~q ),
	.cin(gnd),
	.combout(\Equal9~0_combout ),
	.cout());
defparam \Equal9~0 .lut_mask = 16'h000A;
defparam \Equal9~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal8~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\id_inst[4]~q ),
	.datad(\id_inst[12]~q ),
	.cin(gnd),
	.combout(\Equal8~1_combout ),
	.cout());
defparam \Equal8~1 .lut_mask = 16'h000F;
defparam \Equal8~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal8~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\id_inst[14]~q ),
	.datad(\id_inst[13]~q ),
	.cin(gnd),
	.combout(\Equal8~0_combout ),
	.cout());
defparam \Equal8~0 .lut_mask = 16'h000F;
defparam \Equal8~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal10~0 (
	.dataa(\id_inst[5]~q ),
	.datab(\ex_ctrl_mem_wr~7_combout ),
	.datac(\id_inst[12]~q ),
	.datad(\Equal8~0_combout ),
	.cin(gnd),
	.combout(\Equal10~0_combout ),
	.cout());
defparam \Equal10~0 .lut_mask = 16'h8000;
defparam \Equal10~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal10~1 (
	.dataa(\id_inst[6]~q ),
	.datab(\Equal10~0_combout ),
	.datac(gnd),
	.datad(\id_inst[4]~q ),
	.cin(gnd),
	.combout(\Equal10~1_combout ),
	.cout());
defparam \Equal10~1 .lut_mask = 16'h0088;
defparam \Equal10~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~4 (
	.dataa(\Equal7~0_combout ),
	.datab(\Equal9~0_combout ),
	.datac(\Equal8~1_combout ),
	.datad(\Equal10~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~4_combout ),
	.cout());
defparam \ex_ctrl_alu_func~4 .lut_mask = 16'h007F;
defparam \ex_ctrl_alu_func~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_ctrl_br_type[2]~11 (
	.dataa(\id_inst[12]~q ),
	.datab(\id_inst[13]~q ),
	.datac(\Equal11~0_combout ),
	.datad(\ex_ctrl_alu_func~4_combout ),
	.cin(gnd),
	.combout(\id_ctrl_br_type[2]~11_combout ),
	.cout());
defparam \id_ctrl_br_type[2]~11 .lut_mask = 16'h20FF;
defparam \id_ctrl_br_type[2]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal5~0 (
	.dataa(\id_inst[2]~q ),
	.datab(\id_inst[0]~q ),
	.datac(\id_inst[1]~q ),
	.datad(\id_inst[3]~q ),
	.cin(gnd),
	.combout(\Equal5~0_combout ),
	.cout());
defparam \Equal5~0 .lut_mask = 16'h0080;
defparam \Equal5~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal8~2 (
	.dataa(\Equal5~0_combout ),
	.datab(\Equal7~0_combout ),
	.datac(\Equal8~0_combout ),
	.datad(\Equal8~1_combout ),
	.cin(gnd),
	.combout(\Equal8~2_combout ),
	.cout());
defparam \Equal8~2 .lut_mask = 16'h8000;
defparam \Equal8~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_GEN_15~0 (
	.dataa(\id_inst[12]~q ),
	.datab(\id_inst[13]~q ),
	.datac(gnd),
	.datad(\Equal11~0_combout ),
	.cin(gnd),
	.combout(\_GEN_15~0_combout ),
	.cout());
defparam \_GEN_15~0 .lut_mask = 16'h88FF;
defparam \_GEN_15~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal53~0 (
	.dataa(\id_inst[3]~q ),
	.datab(\id_inst[2]~q ),
	.datac(\id_inst[0]~q ),
	.datad(\id_inst[1]~q ),
	.cin(gnd),
	.combout(\Equal53~0_combout ),
	.cout());
defparam \Equal53~0 .lut_mask = 16'h8000;
defparam \Equal53~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal6~3 (
	.dataa(\id_inst[4]~q ),
	.datab(\id_inst[5]~q ),
	.datac(\id_inst[6]~q ),
	.datad(\Equal5~0_combout ),
	.cin(gnd),
	.combout(\Equal6~3_combout ),
	.cout());
defparam \Equal6~3 .lut_mask = 16'h0200;
defparam \Equal6~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_op1~2 (
	.dataa(\id_inst[4]~q ),
	.datab(\Equal7~0_combout ),
	.datac(\Equal53~0_combout ),
	.datad(\Equal6~3_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_op1~2_combout ),
	.cout());
defparam \ex_ctrl_alu_op1~2 .lut_mask = 16'hFF40;
defparam \ex_ctrl_alu_op1~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal5~1 (
	.dataa(\Equal5~0_combout ),
	.datab(\id_inst[4]~q ),
	.datac(\id_inst[5]~q ),
	.datad(\id_inst[6]~q ),
	.cin(gnd),
	.combout(\Equal5~1_combout ),
	.cout());
defparam \Equal5~1 .lut_mask = 16'h0080;
defparam \Equal5~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_imm_type~14 (
	.dataa(\_GEN_15~0_combout ),
	.datab(\ex_ctrl_alu_func~4_combout ),
	.datac(\ex_ctrl_alu_op1~2_combout ),
	.datad(\Equal5~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_imm_type~14_combout ),
	.cout());
defparam \ex_ctrl_imm_type~14 .lut_mask = 16'h0008;
defparam \ex_ctrl_imm_type~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_ctrl_br_type[0]~4 (
	.dataa(\Equal8~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ex_ctrl_imm_type~14_combout ),
	.cin(gnd),
	.combout(\id_ctrl_br_type[0]~4_combout ),
	.cout());
defparam \id_ctrl_br_type[0]~4 .lut_mask = 16'hAAFF;
defparam \id_ctrl_br_type[0]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_ctrl_br_type[2]~5 (
	.dataa(\Equal14~0_combout ),
	.datab(\id_ctrl_br_type[2]~11_combout ),
	.datac(\id_ctrl_br_type[0]~4_combout ),
	.datad(\Equal5~1_combout ),
	.cin(gnd),
	.combout(\id_ctrl_br_type[2]~5_combout ),
	.cout());
defparam \id_ctrl_br_type[2]~5 .lut_mask = 16'h0ACA;
defparam \id_ctrl_br_type[2]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_br_type~0 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_ctrl_br_type[2]~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_ctrl_br_type~0_combout ),
	.cout());
defparam \ex_ctrl_br_type~0 .lut_mask = 16'h8080;
defparam \ex_ctrl_br_type~0 .sum_lutc_input = "datac";

dffeas \ex_ctrl_br_type[2] (
	.clk(clk_clk),
	.d(\ex_ctrl_br_type~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_br_type[2]~q ),
	.prn(vcc));
defparam \ex_ctrl_br_type[2] .is_wysiwyg = "true";
defparam \ex_ctrl_br_type[2] .power_up = "low";

cyclone10lp_lcell_comb \mem_ctrl_br_type~0 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_ctrl_br_type[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_ctrl_br_type~0_combout ),
	.cout());
defparam \mem_ctrl_br_type~0 .lut_mask = 16'h8888;
defparam \mem_ctrl_br_type~0 .sum_lutc_input = "datac";

dffeas \mem_ctrl_br_type[2] (
	.clk(clk_clk),
	.d(\mem_ctrl_br_type~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_ctrl_br_type[2]~q ),
	.prn(vcc));
defparam \mem_ctrl_br_type[2] .is_wysiwyg = "true";
defparam \mem_ctrl_br_type[2] .power_up = "low";

cyclone10lp_lcell_comb \id_pc[7]~31 (
	.dataa(\inst_kill~0_combout ),
	.datab(\csr|io_expt~combout ),
	.datac(\csr|mcause[0]~6_combout ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\id_pc[7]~31_combout ),
	.cout());
defparam \id_pc[7]~31 .lut_mask = 16'h7FFF;
defparam \id_pc[7]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_br_type~1 (
	.dataa(\id_pc[7]~31_combout ),
	.datab(\Equal11~0_combout ),
	.datac(gnd),
	.datad(\id_inst[12]~q ),
	.cin(gnd),
	.combout(\ex_ctrl_br_type~1_combout ),
	.cout());
defparam \ex_ctrl_br_type~1 .lut_mask = 16'h0044;
defparam \ex_ctrl_br_type~1 .sum_lutc_input = "datac";

dffeas \ex_ctrl_br_type[3] (
	.clk(clk_clk),
	.d(\ex_ctrl_br_type~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_br_type[3]~q ),
	.prn(vcc));
defparam \ex_ctrl_br_type[3] .is_wysiwyg = "true";
defparam \ex_ctrl_br_type[3] .power_up = "low";

cyclone10lp_lcell_comb \mem_ctrl_br_type~1 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_ctrl_br_type[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_ctrl_br_type~1_combout ),
	.cout());
defparam \mem_ctrl_br_type~1 .lut_mask = 16'h8888;
defparam \mem_ctrl_br_type~1 .sum_lutc_input = "datac";

dffeas \mem_ctrl_br_type[3] (
	.clk(clk_clk),
	.d(\mem_ctrl_br_type~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_ctrl_br_type[3]~q ),
	.prn(vcc));
defparam \mem_ctrl_br_type[3] .is_wysiwyg = "true";
defparam \mem_ctrl_br_type[3] .power_up = "low";

cyclone10lp_lcell_comb \Equal2~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\mem_ctrl_br_type[2]~q ),
	.datad(\mem_ctrl_br_type[3]~q ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'h000F;
defparam \Equal2~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~11 (
	.dataa(\id_inst[21]~q ),
	.datab(\_T_1778~combout ),
	.datac(q_a_21),
	.datad(\id_inst~0_combout ),
	.cin(gnd),
	.combout(\id_inst~11_combout ),
	.cout());
defparam \id_inst~11 .lut_mask = 16'hEAC0;
defparam \id_inst~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~12 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\id_inst~11_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~12_combout ),
	.cout());
defparam \id_inst~12 .lut_mask = 16'h8888;
defparam \id_inst~12 .sum_lutc_input = "datac";

dffeas \id_inst[21] (
	.clk(clk_clk),
	.d(\id_inst~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\id_inst[21]~q ),
	.prn(vcc));
defparam \id_inst[21] .is_wysiwyg = "true";
defparam \id_inst[21] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~3 (
	.dataa(\id_inst[15]~q ),
	.datab(\_T_1778~combout ),
	.datac(q_a_15),
	.datad(\id_inst~0_combout ),
	.cin(gnd),
	.combout(\id_inst~3_combout ),
	.cout());
defparam \id_inst~3 .lut_mask = 16'hEAC0;
defparam \id_inst~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~4 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\id_inst~3_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~4_combout ),
	.cout());
defparam \id_inst~4 .lut_mask = 16'h8888;
defparam \id_inst~4 .sum_lutc_input = "datac";

dffeas \id_inst[15] (
	.clk(clk_clk),
	.d(\id_inst~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\id_inst[15]~q ),
	.prn(vcc));
defparam \id_inst[15] .is_wysiwyg = "true";
defparam \id_inst[15] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~1 (
	.dataa(\id_inst[16]~q ),
	.datab(\_T_1778~combout ),
	.datac(q_a_16),
	.datad(\id_inst~0_combout ),
	.cin(gnd),
	.combout(\id_inst~1_combout ),
	.cout());
defparam \id_inst~1 .lut_mask = 16'hEAC0;
defparam \id_inst~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\id_inst~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~2_combout ),
	.cout());
defparam \id_inst~2 .lut_mask = 16'h8888;
defparam \id_inst~2 .sum_lutc_input = "datac";

dffeas \id_inst[16] (
	.clk(clk_clk),
	.d(\id_inst~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\id_inst[16]~q ),
	.prn(vcc));
defparam \id_inst[16] .is_wysiwyg = "true";
defparam \id_inst[16] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~7 (
	.dataa(\id_inst[17]~q ),
	.datab(\_T_1778~combout ),
	.datac(q_a_17),
	.datad(\id_inst~0_combout ),
	.cin(gnd),
	.combout(\id_inst~7_combout ),
	.cout());
defparam \id_inst~7 .lut_mask = 16'hEAC0;
defparam \id_inst~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~8 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\id_inst~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~8_combout ),
	.cout());
defparam \id_inst~8 .lut_mask = 16'h8888;
defparam \id_inst~8 .sum_lutc_input = "datac";

dffeas \id_inst[17] (
	.clk(clk_clk),
	.d(\id_inst~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\id_inst[17]~q ),
	.prn(vcc));
defparam \id_inst[17] .is_wysiwyg = "true";
defparam \id_inst[17] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~5 (
	.dataa(\id_inst[18]~q ),
	.datab(\_T_1778~combout ),
	.datac(q_a_18),
	.datad(\id_inst~0_combout ),
	.cin(gnd),
	.combout(\id_inst~5_combout ),
	.cout());
defparam \id_inst~5 .lut_mask = 16'hEAC0;
defparam \id_inst~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~6 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\id_inst~5_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~6_combout ),
	.cout());
defparam \id_inst~6 .lut_mask = 16'h8888;
defparam \id_inst~6 .sum_lutc_input = "datac";

dffeas \id_inst[18] (
	.clk(clk_clk),
	.d(\id_inst~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\id_inst[18]~q ),
	.prn(vcc));
defparam \id_inst[18] .is_wysiwyg = "true";
defparam \id_inst[18] .power_up = "low";

cyclone10lp_lcell_comb \ex_rs_0[3]~0 (
	.dataa(\id_inst[15]~q ),
	.datab(\id_inst[16]~q ),
	.datac(\id_inst[17]~q ),
	.datad(\id_inst[18]~q ),
	.cin(gnd),
	.combout(\ex_rs_0[3]~0_combout ),
	.cout());
defparam \ex_rs_0[3]~0 .lut_mask = 16'h0001;
defparam \ex_rs_0[3]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~9 (
	.dataa(\id_inst[19]~q ),
	.datab(\_T_1778~combout ),
	.datac(q_a_19),
	.datad(\id_inst~0_combout ),
	.cin(gnd),
	.combout(\id_inst~9_combout ),
	.cout());
defparam \id_inst~9 .lut_mask = 16'hEAC0;
defparam \id_inst~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~10 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\id_inst~9_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~10_combout ),
	.cout());
defparam \id_inst~10 .lut_mask = 16'h8888;
defparam \id_inst~10 .sum_lutc_input = "datac";

dffeas \id_inst[19] (
	.clk(clk_clk),
	.d(\id_inst~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\id_inst[19]~q ),
	.prn(vcc));
defparam \id_inst[19] .is_wysiwyg = "true";
defparam \id_inst[19] .power_up = "low";

cyclone10lp_lcell_comb \ex_rs_0[3]~1 (
	.dataa(\ex_rs_0[3]~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\id_inst[19]~q ),
	.cin(gnd),
	.combout(\ex_rs_0[3]~1_combout ),
	.cout());
defparam \ex_rs_0[3]~1 .lut_mask = 16'h00AA;
defparam \ex_rs_0[3]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~19 (
	.dataa(\id_inst[24]~q ),
	.datab(\_T_1778~combout ),
	.datac(q_a_24),
	.datad(\id_inst~0_combout ),
	.cin(gnd),
	.combout(\id_inst~19_combout ),
	.cout());
defparam \id_inst~19 .lut_mask = 16'hEAC0;
defparam \id_inst~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~20 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\id_inst~19_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~20_combout ),
	.cout());
defparam \id_inst~20 .lut_mask = 16'h8888;
defparam \id_inst~20 .sum_lutc_input = "datac";

dffeas \id_inst[24] (
	.clk(clk_clk),
	.d(\id_inst~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\id_inst[24]~q ),
	.prn(vcc));
defparam \id_inst[24] .is_wysiwyg = "true";
defparam \id_inst[24] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~17 (
	.dataa(\id_inst[22]~q ),
	.datab(\_T_1778~combout ),
	.datac(q_a_22),
	.datad(\id_inst~0_combout ),
	.cin(gnd),
	.combout(\id_inst~17_combout ),
	.cout());
defparam \id_inst~17 .lut_mask = 16'hEAC0;
defparam \id_inst~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~18 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\id_inst~17_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~18_combout ),
	.cout());
defparam \id_inst~18 .lut_mask = 16'h8888;
defparam \id_inst~18 .sum_lutc_input = "datac";

dffeas \id_inst[22] (
	.clk(clk_clk),
	.d(\id_inst~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\id_inst[22]~q ),
	.prn(vcc));
defparam \id_inst[22] .is_wysiwyg = "true";
defparam \id_inst[22] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~15 (
	.dataa(\id_inst[23]~q ),
	.datab(\_T_1778~combout ),
	.datac(q_a_23),
	.datad(\id_inst~0_combout ),
	.cin(gnd),
	.combout(\id_inst~15_combout ),
	.cout());
defparam \id_inst~15 .lut_mask = 16'hEAC0;
defparam \id_inst~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~16 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\id_inst~15_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~16_combout ),
	.cout());
defparam \id_inst~16 .lut_mask = 16'h8888;
defparam \id_inst~16 .sum_lutc_input = "datac";

dffeas \id_inst[23] (
	.clk(clk_clk),
	.d(\id_inst~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\id_inst[23]~q ),
	.prn(vcc));
defparam \id_inst[23] .is_wysiwyg = "true";
defparam \id_inst[23] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~25 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_7),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~25_combout ),
	.cout());
defparam \id_inst~25 .lut_mask = 16'h8080;
defparam \id_inst~25 .sum_lutc_input = "datac";

dffeas \id_inst[7] (
	.clk(clk_clk),
	.d(\id_inst~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[7]~q ),
	.prn(vcc));
defparam \id_inst[7] .is_wysiwyg = "true";
defparam \id_inst[7] .power_up = "low";

cyclone10lp_lcell_comb \Equal48~0 (
	.dataa(\id_inst[24]~q ),
	.datab(\id_inst[22]~q ),
	.datac(\id_inst[23]~q ),
	.datad(\id_inst[7]~q ),
	.cin(gnd),
	.combout(\Equal48~0_combout ),
	.cout());
defparam \Equal48~0 .lut_mask = 16'h0001;
defparam \Equal48~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~26 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_8),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~26_combout ),
	.cout());
defparam \id_inst~26 .lut_mask = 16'h8080;
defparam \id_inst~26 .sum_lutc_input = "datac";

dffeas \id_inst[8] (
	.clk(clk_clk),
	.d(\id_inst~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[8]~q ),
	.prn(vcc));
defparam \id_inst[8] .is_wysiwyg = "true";
defparam \id_inst[8] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~27 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_9),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~27_combout ),
	.cout());
defparam \id_inst~27 .lut_mask = 16'h8080;
defparam \id_inst~27 .sum_lutc_input = "datac";

dffeas \id_inst[9] (
	.clk(clk_clk),
	.d(\id_inst~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[9]~q ),
	.prn(vcc));
defparam \id_inst[9] .is_wysiwyg = "true";
defparam \id_inst[9] .power_up = "low";

cyclone10lp_lcell_comb \Equal48~1 (
	.dataa(\Equal7~0_combout ),
	.datab(\Equal48~0_combout ),
	.datac(\id_inst[8]~q ),
	.datad(\id_inst[9]~q ),
	.cin(gnd),
	.combout(\Equal48~1_combout ),
	.cout());
defparam \Equal48~1 .lut_mask = 16'h0008;
defparam \Equal48~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~29 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_10),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~29_combout ),
	.cout());
defparam \id_inst~29 .lut_mask = 16'h8080;
defparam \id_inst~29 .sum_lutc_input = "datac";

dffeas \id_inst[10] (
	.clk(clk_clk),
	.d(\id_inst~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[10]~q ),
	.prn(vcc));
defparam \id_inst[10] .is_wysiwyg = "true";
defparam \id_inst[10] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~30 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_11),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~30_combout ),
	.cout());
defparam \id_inst~30 .lut_mask = 16'h8080;
defparam \id_inst~30 .sum_lutc_input = "datac";

dffeas \id_inst[11] (
	.clk(clk_clk),
	.d(\id_inst~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[11]~q ),
	.prn(vcc));
defparam \id_inst[11] .is_wysiwyg = "true";
defparam \id_inst[11] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~31 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_25),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~31_combout ),
	.cout());
defparam \id_inst~31 .lut_mask = 16'h8080;
defparam \id_inst~31 .sum_lutc_input = "datac";

dffeas \id_inst[25] (
	.clk(clk_clk),
	.d(\id_inst~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[25]~q ),
	.prn(vcc));
defparam \id_inst[25] .is_wysiwyg = "true";
defparam \id_inst[25] .power_up = "low";

cyclone10lp_lcell_comb \Equal48~2 (
	.dataa(\id_inst[12]~q ),
	.datab(\id_inst[10]~q ),
	.datac(\id_inst[11]~q ),
	.datad(\id_inst[25]~q ),
	.cin(gnd),
	.combout(\Equal48~2_combout ),
	.cout());
defparam \Equal48~2 .lut_mask = 16'h0001;
defparam \Equal48~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~32 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_30),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~32_combout ),
	.cout());
defparam \id_inst~32 .lut_mask = 16'h8080;
defparam \id_inst~32 .sum_lutc_input = "datac";

dffeas \id_inst[30] (
	.clk(clk_clk),
	.d(\id_inst~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[30]~q ),
	.prn(vcc));
defparam \id_inst[30] .is_wysiwyg = "true";
defparam \id_inst[30] .power_up = "low";

cyclone10lp_lcell_comb \Equal48~3 (
	.dataa(\ex_rs_0[3]~1_combout ),
	.datab(\Equal48~1_combout ),
	.datac(\Equal48~2_combout ),
	.datad(\id_inst[30]~q ),
	.cin(gnd),
	.combout(\Equal48~3_combout ),
	.cout());
defparam \Equal48~3 .lut_mask = 16'h0080;
defparam \Equal48~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~38 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_26),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~38_combout ),
	.cout());
defparam \id_inst~38 .lut_mask = 16'h8080;
defparam \id_inst~38 .sum_lutc_input = "datac";

dffeas \id_inst[26] (
	.clk(clk_clk),
	.d(\id_inst~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[26]~q ),
	.prn(vcc));
defparam \id_inst[26] .is_wysiwyg = "true";
defparam \id_inst[26] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~39 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_27),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~39_combout ),
	.cout());
defparam \id_inst~39 .lut_mask = 16'h8080;
defparam \id_inst~39 .sum_lutc_input = "datac";

dffeas \id_inst[27] (
	.clk(clk_clk),
	.d(\id_inst~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[27]~q ),
	.prn(vcc));
defparam \id_inst[27] .is_wysiwyg = "true";
defparam \id_inst[27] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~40 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_31),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~40_combout ),
	.cout());
defparam \id_inst~40 .lut_mask = 16'h8080;
defparam \id_inst~40 .sum_lutc_input = "datac";

dffeas \id_inst[31] (
	.clk(clk_clk),
	.d(\id_inst~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[31]~q ),
	.prn(vcc));
defparam \id_inst[31] .is_wysiwyg = "true";
defparam \id_inst[31] .power_up = "low";

cyclone10lp_lcell_comb \Equal49~0 (
	.dataa(\id_inst[4]~q ),
	.datab(\id_inst[26]~q ),
	.datac(\id_inst[27]~q ),
	.datad(\id_inst[31]~q ),
	.cin(gnd),
	.combout(\Equal49~0_combout ),
	.cout());
defparam \Equal49~0 .lut_mask = 16'h0002;
defparam \Equal49~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~41 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_28),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~41_combout ),
	.cout());
defparam \id_inst~41 .lut_mask = 16'h8080;
defparam \id_inst~41 .sum_lutc_input = "datac";

dffeas \id_inst[28] (
	.clk(clk_clk),
	.d(\id_inst~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[28]~q ),
	.prn(vcc));
defparam \id_inst[28] .is_wysiwyg = "true";
defparam \id_inst[28] .power_up = "low";

cyclone10lp_lcell_comb \id_inst~13 (
	.dataa(\id_inst[20]~q ),
	.datab(\_T_1778~combout ),
	.datac(q_a_20),
	.datad(\id_inst~0_combout ),
	.cin(gnd),
	.combout(\id_inst~13_combout ),
	.cout());
defparam \id_inst~13 .lut_mask = 16'hEAC0;
defparam \id_inst~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~14 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\id_inst~13_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~14_combout ),
	.cout());
defparam \id_inst~14 .lut_mask = 16'h8888;
defparam \id_inst~14 .sum_lutc_input = "datac";

dffeas \id_inst[20] (
	.clk(clk_clk),
	.d(\id_inst~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\id_inst[20]~q ),
	.prn(vcc));
defparam \id_inst[20] .is_wysiwyg = "true";
defparam \id_inst[20] .power_up = "low";

cyclone10lp_lcell_comb \Equal49~1 (
	.dataa(\id_inst[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\id_inst[20]~q ),
	.cin(gnd),
	.combout(\Equal49~1_combout ),
	.cout());
defparam \Equal49~1 .lut_mask = 16'h00AA;
defparam \Equal49~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal49~2 (
	.dataa(\Equal9~0_combout ),
	.datab(\Equal48~3_combout ),
	.datac(\Equal49~0_combout ),
	.datad(\Equal49~1_combout ),
	.cin(gnd),
	.combout(\Equal49~2_combout ),
	.cout());
defparam \Equal49~2 .lut_mask = 16'h8000;
defparam \Equal49~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_inst~42 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(q_a_29),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_inst~42_combout ),
	.cout());
defparam \id_inst~42 .lut_mask = 16'h8080;
defparam \id_inst~42 .sum_lutc_input = "datac";

dffeas \id_inst[29] (
	.clk(clk_clk),
	.d(\id_inst~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_inst[29]~q ),
	.prn(vcc));
defparam \id_inst[29] .is_wysiwyg = "true";
defparam \id_inst[29] .power_up = "low";

cyclone10lp_lcell_comb \Equal49~3 (
	.dataa(\id_inst[21]~q ),
	.datab(\Equal49~2_combout ),
	.datac(\id_inst[29]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal49~3_combout ),
	.cout());
defparam \Equal49~3 .lut_mask = 16'h8080;
defparam \Equal49~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal15~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\id_inst[5]~q ),
	.datad(\id_inst[6]~q ),
	.cin(gnd),
	.combout(\Equal15~0_combout ),
	.cout());
defparam \Equal15~0 .lut_mask = 16'h000F;
defparam \Equal15~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal17~0 (
	.dataa(\ex_ctrl_mem_wr~7_combout ),
	.datab(\id_inst[13]~q ),
	.datac(\Equal15~0_combout ),
	.datad(\id_inst[14]~q ),
	.cin(gnd),
	.combout(\Equal17~0_combout ),
	.cout());
defparam \Equal17~0 .lut_mask = 16'h0080;
defparam \Equal17~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal20~0 (
	.dataa(\id_inst[5]~q ),
	.datab(\Equal9~0_combout ),
	.datac(\Equal8~1_combout ),
	.datad(\id_inst[6]~q ),
	.cin(gnd),
	.combout(\Equal20~0_combout ),
	.cout());
defparam \Equal20~0 .lut_mask = 16'h0080;
defparam \Equal20~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_imm_type~11 (
	.dataa(\id_inst[4]~q ),
	.datab(\id_inst[6]~q ),
	.datac(\Equal10~0_combout ),
	.datad(\Equal20~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_imm_type~11_combout ),
	.cout());
defparam \ex_ctrl_imm_type~11 .lut_mask = 16'h00EF;
defparam \ex_ctrl_imm_type~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal22~0 (
	.dataa(\id_inst[5]~q ),
	.datab(\ex_ctrl_mem_wr~7_combout ),
	.datac(\id_inst[13]~q ),
	.datad(\id_inst[14]~q ),
	.cin(gnd),
	.combout(\Equal22~0_combout ),
	.cout());
defparam \Equal22~0 .lut_mask = 16'h0080;
defparam \Equal22~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_imm_type~12 (
	.dataa(\ex_ctrl_imm_type~11_combout ),
	.datab(\id_inst[6]~q ),
	.datac(\Equal8~1_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_imm_type~12_combout ),
	.cout());
defparam \ex_ctrl_imm_type~12 .lut_mask = 16'h8AAA;
defparam \ex_ctrl_imm_type~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal16~0 (
	.dataa(\id_inst[12]~q ),
	.datab(\id_inst[4]~q ),
	.datac(\id_inst[5]~q ),
	.datad(\id_inst[6]~q ),
	.cin(gnd),
	.combout(\Equal16~0_combout ),
	.cout());
defparam \Equal16~0 .lut_mask = 16'h0002;
defparam \Equal16~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mask_type~1 (
	.dataa(\Equal9~0_combout ),
	.datab(\Equal16~0_combout ),
	.datac(\Equal8~1_combout ),
	.datad(\Equal17~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_mask_type~1_combout ),
	.cout());
defparam \ex_ctrl_mask_type~1 .lut_mask = 16'h0777;
defparam \ex_ctrl_mask_type~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal18~1 (
	.dataa(\id_inst[14]~q ),
	.datab(\ex_ctrl_mem_wr~7_combout ),
	.datac(\Equal15~0_combout ),
	.datad(\id_inst[13]~q ),
	.cin(gnd),
	.combout(\Equal18~1_combout ),
	.cout());
defparam \Equal18~1 .lut_mask = 16'h0080;
defparam \Equal18~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mask_type~2 (
	.dataa(\id_inst[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal18~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_mask_type~2_combout ),
	.cout());
defparam \ex_ctrl_mask_type~2 .lut_mask = 16'hAAFF;
defparam \ex_ctrl_mask_type~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal15~1 (
	.dataa(\ex_ctrl_mem_wr~7_combout ),
	.datab(\Equal8~0_combout ),
	.datac(\Equal8~1_combout ),
	.datad(\Equal15~0_combout ),
	.cin(gnd),
	.combout(\Equal15~1_combout ),
	.cout());
defparam \Equal15~1 .lut_mask = 16'h8000;
defparam \Equal15~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3091~0 (
	.dataa(\ex_ctrl_imm_type~12_combout ),
	.datab(\ex_ctrl_mask_type~1_combout ),
	.datac(\ex_ctrl_mask_type~2_combout ),
	.datad(\Equal15~1_combout ),
	.cin(gnd),
	.combout(\_T_3091~0_combout ),
	.cout());
defparam \_T_3091~0 .lut_mask = 16'h0080;
defparam \_T_3091~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal6~2 (
	.dataa(\id_inst[4]~q ),
	.datab(gnd),
	.datac(\id_inst[5]~q ),
	.datad(\id_inst[6]~q ),
	.cin(gnd),
	.combout(\Equal6~2_combout ),
	.cout());
defparam \Equal6~2 .lut_mask = 16'h000A;
defparam \Equal6~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~9 (
	.dataa(\_T_3091~0_combout ),
	.datab(\id_inst[12]~q ),
	.datac(\Equal9~0_combout ),
	.datad(\Equal6~2_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~9_combout ),
	.cout());
defparam \ex_ctrl_alu_func~9 .lut_mask = 16'h8AAA;
defparam \ex_ctrl_alu_func~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_2062[1]~0 (
	.dataa(\id_inst[4]~q ),
	.datab(\Equal17~0_combout ),
	.datac(\id_inst[12]~q ),
	.datad(\ex_ctrl_alu_func~9_combout ),
	.cin(gnd),
	.combout(\_T_2062[1]~0_combout ),
	.cout());
defparam \_T_2062[1]~0 .lut_mask = 16'h08FF;
defparam \_T_2062[1]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_ctrl_br_type[1]~6 (
	.dataa(\Equal14~0_combout ),
	.datab(\Equal49~3_combout ),
	.datac(\_T_2062[1]~0_combout ),
	.datad(\id_ctrl_br_type[0]~4_combout ),
	.cin(gnd),
	.combout(\id_ctrl_br_type[1]~6_combout ),
	.cout());
defparam \id_ctrl_br_type[1]~6 .lut_mask = 16'h00AE;
defparam \id_ctrl_br_type[1]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_ctrl_br_type[1]~12 (
	.dataa(\id_inst[12]~q ),
	.datab(\id_inst[13]~q ),
	.datac(\Equal11~0_combout ),
	.datad(\Equal8~2_combout ),
	.cin(gnd),
	.combout(\id_ctrl_br_type[1]~12_combout ),
	.cout());
defparam \id_ctrl_br_type[1]~12 .lut_mask = 16'h00DF;
defparam \id_ctrl_br_type[1]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_ctrl_br_type[1]~10 (
	.dataa(\id_ctrl_br_type[1]~6_combout ),
	.datab(\id_ctrl_br_type[0]~4_combout ),
	.datac(\Equal5~1_combout ),
	.datad(\id_ctrl_br_type[1]~12_combout ),
	.cin(gnd),
	.combout(\id_ctrl_br_type[1]~10_combout ),
	.cout());
defparam \id_ctrl_br_type[1]~10 .lut_mask = 16'hAAAE;
defparam \id_ctrl_br_type[1]~10 .sum_lutc_input = "datac";

dffeas \ex_ctrl_br_type[1] (
	.clk(clk_clk),
	.d(\id_ctrl_br_type[1]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\id_pc[7]~31_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_br_type[1]~q ),
	.prn(vcc));
defparam \ex_ctrl_br_type[1] .is_wysiwyg = "true";
defparam \ex_ctrl_br_type[1] .power_up = "low";

cyclone10lp_lcell_comb \mem_ctrl_br_type~3 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_ctrl_br_type[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_ctrl_br_type~3_combout ),
	.cout());
defparam \mem_ctrl_br_type~3 .lut_mask = 16'h8888;
defparam \mem_ctrl_br_type~3 .sum_lutc_input = "datac";

dffeas \mem_ctrl_br_type[1] (
	.clk(clk_clk),
	.d(\mem_ctrl_br_type~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_ctrl_br_type[1]~q ),
	.prn(vcc));
defparam \mem_ctrl_br_type[1] .is_wysiwyg = "true";
defparam \mem_ctrl_br_type[1] .power_up = "low";

cyclone10lp_lcell_comb \inst_kill~1 (
	.dataa(\inst_kill~0_combout ),
	.datab(\csr|io_expt~0_combout ),
	.datac(gnd),
	.datad(\csr|isEcall~0_combout ),
	.cin(gnd),
	.combout(\inst_kill~1_combout ),
	.cout());
defparam \inst_kill~1 .lut_mask = 16'h0088;
defparam \inst_kill~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal9~1 (
	.dataa(\ex_ctrl_mem_wr~7_combout ),
	.datab(\Equal8~0_combout ),
	.datac(\id_inst[4]~q ),
	.datad(\id_inst[12]~q ),
	.cin(gnd),
	.combout(\Equal9~1_combout ),
	.cout());
defparam \Equal9~1 .lut_mask = 16'h0008;
defparam \Equal9~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~10 (
	.dataa(\ex_ctrl_alu_op1~2_combout ),
	.datab(\Equal7~0_combout ),
	.datac(\Equal9~1_combout ),
	.datad(\Equal8~2_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~10_combout ),
	.cout());
defparam \ex_ctrl_alu_func~10 .lut_mask = 16'h0015;
defparam \ex_ctrl_alu_func~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal26~0 (
	.dataa(\id_inst[4]~q ),
	.datab(\Equal18~1_combout ),
	.datac(gnd),
	.datad(\id_inst[12]~q ),
	.cin(gnd),
	.combout(\Equal26~0_combout ),
	.cout());
defparam \Equal26~0 .lut_mask = 16'h0088;
defparam \Equal26~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal13~0 (
	.dataa(\id_inst[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\id_inst[12]~q ),
	.cin(gnd),
	.combout(\Equal13~0_combout ),
	.cout());
defparam \Equal13~0 .lut_mask = 16'h00AA;
defparam \Equal13~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal27~0 (
	.dataa(\id_inst[14]~q ),
	.datab(\ex_ctrl_mem_wr~7_combout ),
	.datac(\Equal13~0_combout ),
	.datad(\Equal6~2_combout ),
	.cin(gnd),
	.combout(\Equal27~0_combout ),
	.cout());
defparam \Equal27~0 .lut_mask = 16'h8000;
defparam \Equal27~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~34 (
	.dataa(\id_inst[4]~q ),
	.datab(\Equal17~0_combout ),
	.datac(\Equal26~0_combout ),
	.datad(\Equal27~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~34_combout ),
	.cout());
defparam \ex_ctrl_alu_func~34 .lut_mask = 16'h0007;
defparam \ex_ctrl_alu_func~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal28~0 (
	.dataa(\id_inst[4]~q ),
	.datab(\id_inst[12]~q ),
	.datac(\id_inst[5]~q ),
	.datad(\id_inst[6]~q ),
	.cin(gnd),
	.combout(\Equal28~0_combout ),
	.cout());
defparam \Equal28~0 .lut_mask = 16'h0008;
defparam \Equal28~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal28~1 (
	.dataa(\id_inst[14]~q ),
	.datab(\ex_ctrl_mem_wr~7_combout ),
	.datac(\id_inst[13]~q ),
	.datad(\Equal28~0_combout ),
	.cin(gnd),
	.combout(\Equal28~1_combout ),
	.cout());
defparam \Equal28~1 .lut_mask = 16'h8000;
defparam \Equal28~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal12~0 (
	.dataa(\id_inst[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\id_inst[13]~q ),
	.cin(gnd),
	.combout(\Equal12~0_combout ),
	.cout());
defparam \Equal12~0 .lut_mask = 16'h00AA;
defparam \Equal12~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal29~0 (
	.dataa(\ex_ctrl_mem_wr~7_combout ),
	.datab(\Equal49~0_combout ),
	.datac(\id_inst[28]~q ),
	.datad(\id_inst[29]~q ),
	.cin(gnd),
	.combout(\Equal29~0_combout ),
	.cout());
defparam \Equal29~0 .lut_mask = 16'h0008;
defparam \Equal29~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal32~0 (
	.dataa(\id_inst[5]~q ),
	.datab(\Equal29~0_combout ),
	.datac(\id_inst[6]~q ),
	.datad(\id_inst[25]~q ),
	.cin(gnd),
	.combout(\Equal32~0_combout ),
	.cout());
defparam \Equal32~0 .lut_mask = 16'h0008;
defparam \Equal32~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal39~0 (
	.dataa(\id_inst[14]~q ),
	.datab(\Equal12~0_combout ),
	.datac(\id_inst[30]~q ),
	.datad(\Equal32~0_combout ),
	.cin(gnd),
	.combout(\Equal39~0_combout ),
	.cout());
defparam \Equal39~0 .lut_mask = 16'h8000;
defparam \Equal39~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal34~0 (
	.dataa(\Equal12~0_combout ),
	.datab(\Equal32~0_combout ),
	.datac(\id_inst[14]~q ),
	.datad(\id_inst[30]~q ),
	.cin(gnd),
	.combout(\Equal34~0_combout ),
	.cout());
defparam \Equal34~0 .lut_mask = 16'h0008;
defparam \Equal34~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal37~0 (
	.dataa(\id_inst[14]~q ),
	.datab(\Equal32~0_combout ),
	.datac(gnd),
	.datad(\id_inst[30]~q ),
	.cin(gnd),
	.combout(\Equal37~0_combout ),
	.cout());
defparam \Equal37~0 .lut_mask = 16'h0088;
defparam \Equal37~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~11 (
	.dataa(\Equal34~0_combout ),
	.datab(\id_inst[12]~q ),
	.datac(\Equal37~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~11_combout ),
	.cout());
defparam \ex_ctrl_alu_func~11 .lut_mask = 16'hEAEA;
defparam \ex_ctrl_alu_func~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal18~0 (
	.dataa(gnd),
	.datab(\id_inst[5]~q ),
	.datac(\id_inst[6]~q ),
	.datad(\id_inst[13]~q ),
	.cin(gnd),
	.combout(\Equal18~0_combout ),
	.cout());
defparam \Equal18~0 .lut_mask = 16'h0003;
defparam \Equal18~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal29~1 (
	.dataa(\id_inst[12]~q ),
	.datab(\Equal18~0_combout ),
	.datac(\Equal29~0_combout ),
	.datad(\id_inst[30]~q ),
	.cin(gnd),
	.combout(\Equal29~1_combout ),
	.cout());
defparam \Equal29~1 .lut_mask = 16'h0080;
defparam \Equal29~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal31~0 (
	.dataa(\id_inst[30]~q ),
	.datab(\Equal29~0_combout ),
	.datac(\id_inst[6]~q ),
	.datad(\id_inst[13]~q ),
	.cin(gnd),
	.combout(\Equal31~0_combout ),
	.cout());
defparam \Equal31~0 .lut_mask = 16'h0008;
defparam \Equal31~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal31~1 (
	.dataa(\id_inst[14]~q ),
	.datab(\id_inst[12]~q ),
	.datac(\Equal31~0_combout ),
	.datad(\id_inst[5]~q ),
	.cin(gnd),
	.combout(\Equal31~1_combout ),
	.cout());
defparam \Equal31~1 .lut_mask = 16'h0080;
defparam \Equal31~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_op2~5 (
	.dataa(\id_inst[25]~q ),
	.datab(\id_inst[14]~q ),
	.datac(\Equal29~1_combout ),
	.datad(\Equal31~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_op2~5_combout ),
	.cout());
defparam \ex_ctrl_alu_op2~5 .lut_mask = 16'h002F;
defparam \ex_ctrl_alu_op2~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~12 (
	.dataa(\Equal28~1_combout ),
	.datab(\Equal39~0_combout ),
	.datac(\ex_ctrl_alu_func~11_combout ),
	.datad(\ex_ctrl_alu_op2~5_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~12_combout ),
	.cout());
defparam \ex_ctrl_alu_func~12 .lut_mask = 16'hFEFF;
defparam \ex_ctrl_alu_func~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~13 (
	.dataa(\Equal14~0_combout ),
	.datab(\ex_ctrl_alu_func~9_combout ),
	.datac(\ex_ctrl_alu_func~34_combout ),
	.datad(\ex_ctrl_alu_func~12_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~13_combout ),
	.cout());
defparam \ex_ctrl_alu_func~13 .lut_mask = 16'hEAAA;
defparam \ex_ctrl_alu_func~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~14 (
	.dataa(\ex_ctrl_alu_func~13_combout ),
	.datab(\id_inst[12]~q ),
	.datac(\Equal11~0_combout ),
	.datad(\id_inst[13]~q ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~14_combout ),
	.cout());
defparam \ex_ctrl_alu_func~14 .lut_mask = 16'h8ACA;
defparam \ex_ctrl_alu_func~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~15 (
	.dataa(\Equal5~1_combout ),
	.datab(\ex_ctrl_alu_func~10_combout ),
	.datac(\Equal10~1_combout ),
	.datad(\ex_ctrl_alu_func~14_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~15_combout ),
	.cout());
defparam \ex_ctrl_alu_func~15 .lut_mask = 16'hEEEA;
defparam \ex_ctrl_alu_func~15 .sum_lutc_input = "datac";

dffeas \ex_ctrl_alu_func[0] (
	.clk(clk_clk),
	.d(\ex_ctrl_alu_func~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\id_pc[7]~31_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_alu_func[0]~q ),
	.prn(vcc));
defparam \ex_ctrl_alu_func[0] .is_wysiwyg = "true";
defparam \ex_ctrl_alu_func[0] .power_up = "low";

cyclone10lp_lcell_comb _GEN_53(
	.dataa(\inst_kill~1_combout ),
	.datab(gnd),
	.datac(\ex_ctrl_alu_func[0]~q ),
	.datad(\alu|_T_125~20_combout ),
	.cin(gnd),
	.combout(\_GEN_53~combout ),
	.cout());
defparam _GEN_53.lut_mask = 16'h0AA0;
defparam _GEN_53.sum_lutc_input = "datac";

dffeas mem_alu_cmp_out(
	.clk(clk_clk),
	.d(\_GEN_53~combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_cmp_out~q ),
	.prn(vcc));
defparam mem_alu_cmp_out.is_wysiwyg = "true";
defparam mem_alu_cmp_out.power_up = "low";

cyclone10lp_lcell_comb \inst_kill~0 (
	.dataa(\Equal2~0_combout ),
	.datab(\mem_ctrl_br_type[0]~q ),
	.datac(\mem_ctrl_br_type[1]~q ),
	.datad(\mem_alu_cmp_out~q ),
	.cin(gnd),
	.combout(\inst_kill~0_combout ),
	.cout());
defparam \inst_kill~0 .lut_mask = 16'h0257;
defparam \inst_kill~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_ctrl_mem_wr~7 (
	.dataa(\inst_kill~0_combout ),
	.datab(\csr|io_expt~0_combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(\csr|isEcall~0_combout ),
	.cin(gnd),
	.combout(\mem_ctrl_mem_wr~7_combout ),
	.cout());
defparam \mem_ctrl_mem_wr~7 .lut_mask = 16'h0080;
defparam \mem_ctrl_mem_wr~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_ctrl_br_type[0]~7 (
	.dataa(\id_inst[13]~q ),
	.datab(gnd),
	.datac(\Equal11~0_combout ),
	.datad(\Equal8~2_combout ),
	.cin(gnd),
	.combout(\id_ctrl_br_type[0]~7_combout ),
	.cout());
defparam \id_ctrl_br_type[0]~7 .lut_mask = 16'h00AF;
defparam \id_ctrl_br_type[0]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_ctrl_br_type[0]~8 (
	.dataa(\id_ctrl_br_type[0]~7_combout ),
	.datab(gnd),
	.datac(\Equal10~1_combout ),
	.datad(\Equal6~3_combout ),
	.cin(gnd),
	.combout(\id_ctrl_br_type[0]~8_combout ),
	.cout());
defparam \id_ctrl_br_type[0]~8 .lut_mask = 16'h000A;
defparam \id_ctrl_br_type[0]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \id_ctrl_br_type[0]~9 (
	.dataa(\id_ctrl_br_type[1]~6_combout ),
	.datab(\id_ctrl_br_type[0]~4_combout ),
	.datac(\id_ctrl_br_type[0]~8_combout ),
	.datad(\Equal5~1_combout ),
	.cin(gnd),
	.combout(\id_ctrl_br_type[0]~9_combout ),
	.cout());
defparam \id_ctrl_br_type[0]~9 .lut_mask = 16'hAAEA;
defparam \id_ctrl_br_type[0]~9 .sum_lutc_input = "datac";

dffeas \ex_ctrl_br_type[0] (
	.clk(clk_clk),
	.d(\id_ctrl_br_type[0]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\id_pc[7]~31_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_br_type[0]~q ),
	.prn(vcc));
defparam \ex_ctrl_br_type[0] .is_wysiwyg = "true";
defparam \ex_ctrl_br_type[0] .power_up = "low";

cyclone10lp_lcell_comb \mem_ctrl_br_type~2 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_ctrl_br_type[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_ctrl_br_type~2_combout ),
	.cout());
defparam \mem_ctrl_br_type~2 .lut_mask = 16'h8888;
defparam \mem_ctrl_br_type~2 .sum_lutc_input = "datac";

dffeas \mem_ctrl_br_type[0] (
	.clk(clk_clk),
	.d(\mem_ctrl_br_type~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_ctrl_br_type[0]~q ),
	.prn(vcc));
defparam \mem_ctrl_br_type[0] .is_wysiwyg = "true";
defparam \mem_ctrl_br_type[0] .power_up = "low";

cyclone10lp_lcell_comb \Equal4~0 (
	.dataa(\mem_ctrl_br_type[0]~q ),
	.datab(\mem_ctrl_br_type[1]~q ),
	.datac(\mem_ctrl_br_type[2]~q ),
	.datad(\mem_ctrl_br_type[3]~q ),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
defparam \Equal4~0 .lut_mask = 16'h0008;
defparam \Equal4~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr[0]~0 (
	.dataa(\Equal4~0_combout ),
	.datab(\csr|isEcall~0_combout ),
	.datac(gnd),
	.datad(\csr|io_expt~0_combout ),
	.cin(gnd),
	.combout(\pc_cntr[0]~0_combout ),
	.cout());
defparam \pc_cntr[0]~0 .lut_mask = 16'hEEFF;
defparam \pc_cntr[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_inst~6 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~6_combout ),
	.cout());
defparam \ex_inst~6 .lut_mask = 16'h8080;
defparam \ex_inst~6 .sum_lutc_input = "datac";

dffeas \ex_inst[7] (
	.clk(clk_clk),
	.d(\ex_inst~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[7]~q ),
	.prn(vcc));
defparam \ex_inst[7] .is_wysiwyg = "true";
defparam \ex_inst[7] .power_up = "low";

cyclone10lp_lcell_comb \ex_inst~0 (
	.dataa(\id_inst[15]~q ),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~0_combout ),
	.cout());
defparam \ex_inst~0 .lut_mask = 16'h8080;
defparam \ex_inst~0 .sum_lutc_input = "datac";

dffeas \ex_inst[15] (
	.clk(clk_clk),
	.d(\ex_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[15]~q ),
	.prn(vcc));
defparam \ex_inst[15] .is_wysiwyg = "true";
defparam \ex_inst[15] .power_up = "low";

cyclone10lp_lcell_comb \ex_ctrl_mask_type~0 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(\Equal5~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_mask_type~0_combout ),
	.cout());
defparam \ex_ctrl_mask_type~0 .lut_mask = 16'h0088;
defparam \ex_ctrl_mask_type~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\id_inst[4]~q ),
	.datad(\Equal17~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~6_combout ),
	.cout());
defparam \ex_ctrl_alu_func~6 .lut_mask = 16'h0FFF;
defparam \ex_ctrl_alu_func~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~7 (
	.dataa(\ex_ctrl_alu_func~6_combout ),
	.datab(\Equal28~1_combout ),
	.datac(\Equal26~0_combout ),
	.datad(\Equal27~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~7_combout ),
	.cout());
defparam \ex_ctrl_alu_func~7 .lut_mask = 16'h0002;
defparam \ex_ctrl_alu_func~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3083~0 (
	.dataa(\ex_ctrl_alu_func~7_combout ),
	.datab(\id_inst[12]~q ),
	.datac(\Equal9~0_combout ),
	.datad(\Equal6~2_combout ),
	.cin(gnd),
	.combout(\_T_3083~0_combout ),
	.cout());
defparam \_T_3083~0 .lut_mask = 16'h8AAA;
defparam \_T_3083~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~33 (
	.dataa(\id_inst[4]~q ),
	.datab(\Equal18~1_combout ),
	.datac(\ex_ctrl_mask_type~1_combout ),
	.datad(\Equal15~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~33_combout ),
	.cout());
defparam \ex_ctrl_alu_func~33 .lut_mask = 16'h00B0;
defparam \ex_ctrl_alu_func~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_GEN_15~1 (
	.dataa(\Equal11~0_combout ),
	.datab(\id_inst[12]~q ),
	.datac(\id_inst[13]~q ),
	.datad(\Equal8~2_combout ),
	.cin(gnd),
	.combout(\_GEN_15~1_combout ),
	.cout());
defparam \_GEN_15~1 .lut_mask = 16'h007F;
defparam \_GEN_15~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_GEN_15~2 (
	.dataa(\_GEN_15~0_combout ),
	.datab(\ex_ctrl_alu_func~4_combout ),
	.datac(\ex_ctrl_alu_op1~2_combout ),
	.datad(\_GEN_15~1_combout ),
	.cin(gnd),
	.combout(\_GEN_15~2_combout ),
	.cout());
defparam \_GEN_15~2 .lut_mask = 16'h0800;
defparam \_GEN_15~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_csr_cmd~9 (
	.dataa(\ex_ctrl_imm_type~12_combout ),
	.datab(\ex_ctrl_alu_func~33_combout ),
	.datac(\_GEN_15~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_ctrl_csr_cmd~9_combout ),
	.cout());
defparam \ex_ctrl_csr_cmd~9 .lut_mask = 16'h8080;
defparam \ex_ctrl_csr_cmd~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal43~0 (
	.dataa(\id_inst[4]~q ),
	.datab(\id_inst[14]~q ),
	.datac(\ex_ctrl_mem_wr~7_combout ),
	.datad(\Equal7~0_combout ),
	.cin(gnd),
	.combout(\Equal43~0_combout ),
	.cout());
defparam \Equal43~0 .lut_mask = 16'h8000;
defparam \Equal43~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_imm_type~13 (
	.dataa(gnd),
	.datab(\id_inst[12]~q ),
	.datac(\id_inst[13]~q ),
	.datad(\Equal43~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_imm_type~13_combout ),
	.cout());
defparam \ex_ctrl_imm_type~13 .lut_mask = 16'h03FF;
defparam \ex_ctrl_imm_type~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_imm_type~17 (
	.dataa(\ex_ctrl_mask_type~0_combout ),
	.datab(\_T_3083~0_combout ),
	.datac(\ex_ctrl_csr_cmd~9_combout ),
	.datad(\ex_ctrl_imm_type~13_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_imm_type~17_combout ),
	.cout());
defparam \ex_ctrl_imm_type~17 .lut_mask = 16'h0080;
defparam \ex_ctrl_imm_type~17 .sum_lutc_input = "datac";

dffeas \ex_ctrl_imm_type.101 (
	.clk(clk_clk),
	.d(\ex_ctrl_imm_type~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_imm_type.101~q ),
	.prn(vcc));
defparam \ex_ctrl_imm_type.101 .is_wysiwyg = "true";
defparam \ex_ctrl_imm_type.101 .power_up = "low";

cyclone10lp_lcell_comb \ex_csr_addr~0 (
	.dataa(\id_inst[20]~q ),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_csr_addr~0_combout ),
	.cout());
defparam \ex_csr_addr~0 .lut_mask = 16'h8080;
defparam \ex_csr_addr~0 .sum_lutc_input = "datac";

dffeas \ex_csr_addr[0] (
	.clk(clk_clk),
	.d(\ex_csr_addr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_addr[0]~q ),
	.prn(vcc));
defparam \ex_csr_addr[0] .is_wysiwyg = "true";
defparam \ex_csr_addr[0] .power_up = "low";

cyclone10lp_lcell_comb \ex_ctrl_imm_type~18 (
	.dataa(\ex_ctrl_imm_type~14_combout ),
	.datab(\ex_ctrl_imm_type~12_combout ),
	.datac(gnd),
	.datad(\Equal14~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_imm_type~18_combout ),
	.cout());
defparam \ex_ctrl_imm_type~18 .lut_mask = 16'h0088;
defparam \ex_ctrl_imm_type~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_imm_type~19 (
	.dataa(\Equal8~2_combout ),
	.datab(\ex_ctrl_imm_type~18_combout ),
	.datac(\id_pc[7]~31_combout ),
	.datad(\ex_ctrl_alu_func~33_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_imm_type~19_combout ),
	.cout());
defparam \ex_ctrl_imm_type~19 .lut_mask = 16'hFEFF;
defparam \ex_ctrl_imm_type~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_csr_cmd~10 (
	.dataa(\id_inst[13]~q ),
	.datab(\Equal32~0_combout ),
	.datac(\id_inst[30]~q ),
	.datad(\id_inst[14]~q ),
	.cin(gnd),
	.combout(\ex_csr_cmd~10_combout ),
	.cout());
defparam \ex_csr_cmd~10 .lut_mask = 16'hF3F7;
defparam \ex_csr_cmd~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal32~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\id_inst[14]~q ),
	.datad(\id_inst[12]~q ),
	.cin(gnd),
	.combout(\Equal32~1_combout ),
	.cout());
defparam \Equal32~1 .lut_mask = 16'h000F;
defparam \Equal32~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal33~0 (
	.dataa(\id_inst[5]~q ),
	.datab(\Equal31~0_combout ),
	.datac(\Equal32~1_combout ),
	.datad(\id_inst[25]~q ),
	.cin(gnd),
	.combout(\Equal33~0_combout ),
	.cout());
defparam \Equal33~0 .lut_mask = 16'h0080;
defparam \Equal33~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\Equal33~0_combout ),
	.datad(\Equal39~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~8_combout ),
	.cout());
defparam \ex_ctrl_alu_func~8 .lut_mask = 16'h000F;
defparam \ex_ctrl_alu_func~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal32~2 (
	.dataa(\Equal32~0_combout ),
	.datab(\Equal32~1_combout ),
	.datac(\id_inst[13]~q ),
	.datad(\id_inst[30]~q ),
	.cin(gnd),
	.combout(\Equal32~2_combout ),
	.cout());
defparam \Equal32~2 .lut_mask = 16'h0008;
defparam \Equal32~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_csr_cmd~10 (
	.dataa(\ex_csr_cmd~10_combout ),
	.datab(\ex_ctrl_alu_func~8_combout ),
	.datac(\Equal32~2_combout ),
	.datad(\Equal34~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_csr_cmd~10_combout ),
	.cout());
defparam \ex_ctrl_csr_cmd~10 .lut_mask = 16'h0008;
defparam \ex_ctrl_csr_cmd~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_csr_cmd~14 (
	.dataa(\ex_ctrl_alu_op2~5_combout ),
	.datab(\_T_3083~0_combout ),
	.datac(\ex_ctrl_csr_cmd~9_combout ),
	.datad(\ex_ctrl_csr_cmd~10_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_csr_cmd~14_combout ),
	.cout());
defparam \ex_ctrl_csr_cmd~14 .lut_mask = 16'h7FFF;
defparam \ex_ctrl_csr_cmd~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_imm_type~20 (
	.dataa(\ex_ctrl_imm_type~19_combout ),
	.datab(\ex_ctrl_imm_type~13_combout ),
	.datac(\ex_ctrl_mask_type~0_combout ),
	.datad(\ex_ctrl_csr_cmd~14_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_imm_type~20_combout ),
	.cout());
defparam \ex_ctrl_imm_type~20 .lut_mask = 16'h5535;
defparam \ex_ctrl_imm_type~20 .sum_lutc_input = "datac";

dffeas \ex_ctrl_imm_type.000 (
	.clk(clk_clk),
	.d(\ex_ctrl_imm_type~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_imm_type.000~q ),
	.prn(vcc));
defparam \ex_ctrl_imm_type.000 .is_wysiwyg = "true";
defparam \ex_ctrl_imm_type.000 .power_up = "low";

cyclone10lp_lcell_comb \io_sw_r_ex_imm[0]~2 (
	.dataa(\ex_inst[15]~q ),
	.datab(\ex_ctrl_imm_type.101~q ),
	.datac(\ex_csr_addr[0]~q ),
	.datad(\ex_ctrl_imm_type.000~q ),
	.cin(gnd),
	.combout(\io_sw_r_ex_imm[0]~2_combout ),
	.cout());
defparam \io_sw_r_ex_imm[0]~2 .lut_mask = 16'h88F0;
defparam \io_sw_r_ex_imm[0]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_csr_cmd~5 (
	.dataa(\ex_ctrl_imm_type~11_combout ),
	.datab(\ex_ctrl_alu_func~33_combout ),
	.datac(\_GEN_15~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_csr_cmd~5_combout ),
	.cout());
defparam \ex_csr_cmd~5 .lut_mask = 16'h8080;
defparam \ex_csr_cmd~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mem_wr~8 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\ex_csr_cmd~5_combout ),
	.datad(\Equal5~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_mem_wr~8_combout ),
	.cout());
defparam \ex_ctrl_mem_wr~8 .lut_mask = 16'h0080;
defparam \ex_ctrl_mem_wr~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mem_wr~9 (
	.dataa(\Equal8~1_combout ),
	.datab(\Equal22~0_combout ),
	.datac(\ex_ctrl_mem_wr~8_combout ),
	.datad(\id_inst[6]~q ),
	.cin(gnd),
	.combout(\ex_ctrl_mem_wr~9_combout ),
	.cout());
defparam \ex_ctrl_mem_wr~9 .lut_mask = 16'h0080;
defparam \ex_ctrl_mem_wr~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mask_type~3 (
	.dataa(\ex_ctrl_alu_func~33_combout ),
	.datab(\_GEN_15~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_ctrl_mask_type~3_combout ),
	.cout());
defparam \ex_ctrl_mask_type~3 .lut_mask = 16'h8888;
defparam \ex_ctrl_mask_type~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mem_wr~10 (
	.dataa(\ex_ctrl_mem_wr~9_combout ),
	.datab(\ex_ctrl_mask_type~0_combout ),
	.datac(\ex_ctrl_mask_type~3_combout ),
	.datad(\ex_ctrl_mem_wr~8_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_mem_wr~10_combout ),
	.cout());
defparam \ex_ctrl_mem_wr~10 .lut_mask = 16'hAAEA;
defparam \ex_ctrl_mem_wr~10 .sum_lutc_input = "datac";

dffeas \ex_ctrl_imm_type.001 (
	.clk(clk_clk),
	.d(\ex_ctrl_mem_wr~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_imm_type.001~q ),
	.prn(vcc));
defparam \ex_ctrl_imm_type.001 .is_wysiwyg = "true";
defparam \ex_ctrl_imm_type.001 .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~46 (
	.dataa(\ex_inst[7]~q ),
	.datab(\io_sw_r_ex_imm[0]~2_combout ),
	.datac(\ex_ctrl_imm_type.001~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_imm~46_combout ),
	.cout());
defparam \mem_imm~46 .lut_mask = 16'hAC00;
defparam \mem_imm~46 .sum_lutc_input = "datac";

dffeas \mem_imm[0] (
	.clk(clk_clk),
	.d(\mem_imm~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[0]~q ),
	.prn(vcc));
defparam \mem_imm[0] .is_wysiwyg = "true";
defparam \mem_imm[0] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[0]~0 (
	.dataa(gnd),
	.datab(\mem_imm[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\_T_3862[0]~0_combout ),
	.cout());
defparam \_T_3862[0]~0 .lut_mask = 16'hCCCC;
defparam \_T_3862[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr[0]~1 (
	.dataa(\mem_alu_cmp_out~q ),
	.datab(\Equal2~0_combout ),
	.datac(\Equal4~0_combout ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr[0]~1_combout ),
	.cout());
defparam \pc_cntr[0]~1 .lut_mask = 16'h02FF;
defparam \pc_cntr[0]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~2 (
	.dataa(\pc_cntr[0]~0_combout ),
	.datab(\_T_3862[0]~0_combout ),
	.datac(\pc_cntr[0]~1_combout ),
	.datad(mem_alu_out_0),
	.cin(gnd),
	.combout(\pc_cntr~2_combout ),
	.cout());
defparam \pc_cntr~2 .lut_mask = 16'hE5E0;
defparam \pc_cntr~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~3 (
	.dataa(\csr|mepc[0]~q ),
	.datab(\pc_cntr[0]~0_combout ),
	.datac(\pc_cntr~2_combout ),
	.datad(\csr|mtvec[0]~q ),
	.cin(gnd),
	.combout(\pc_cntr~3_combout ),
	.cout());
defparam \pc_cntr~3 .lut_mask = 16'hF838;
defparam \pc_cntr~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr[0]~4 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\inst_kill~1_combout ),
	.datac(gnd),
	.datad(\csr|mcause[0]~6_combout ),
	.cin(gnd),
	.combout(\pc_cntr[0]~4_combout ),
	.cout());
defparam \pc_cntr[0]~4 .lut_mask = 16'h7755;
defparam \pc_cntr[0]~4 .sum_lutc_input = "datac";

dffeas \pc_cntr[0] (
	.clk(clk_clk),
	.d(\pc_cntr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(\pc_cntr[0]~4_combout ),
	.q(\pc_cntr[0]~q ),
	.prn(vcc));
defparam \pc_cntr[0] .is_wysiwyg = "true";
defparam \pc_cntr[0] .power_up = "low";

cyclone10lp_lcell_comb \id_npc~0 (
	.dataa(\pc_cntr[0]~q ),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~0_combout ),
	.cout());
defparam \id_npc~0 .lut_mask = 16'h8080;
defparam \id_npc~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_inst~5 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[8]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~5_combout ),
	.cout());
defparam \ex_inst~5 .lut_mask = 16'h8080;
defparam \ex_inst~5 .sum_lutc_input = "datac";

dffeas \ex_inst[8] (
	.clk(clk_clk),
	.d(\ex_inst~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[8]~q ),
	.prn(vcc));
defparam \ex_inst[8] .is_wysiwyg = "true";
defparam \ex_inst[8] .power_up = "low";

cyclone10lp_lcell_comb \ex_inst~1 (
	.dataa(\id_inst[16]~q ),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~1_combout ),
	.cout());
defparam \ex_inst~1 .lut_mask = 16'h8080;
defparam \ex_inst~1 .sum_lutc_input = "datac";

dffeas \ex_inst[16] (
	.clk(clk_clk),
	.d(\ex_inst~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[16]~q ),
	.prn(vcc));
defparam \ex_inst[16] .is_wysiwyg = "true";
defparam \ex_inst[16] .power_up = "low";

cyclone10lp_lcell_comb \ex_csr_addr~1 (
	.dataa(\id_inst[21]~q ),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_csr_addr~1_combout ),
	.cout());
defparam \ex_csr_addr~1 .lut_mask = 16'h8080;
defparam \ex_csr_addr~1 .sum_lutc_input = "datac";

dffeas \ex_csr_addr[1] (
	.clk(clk_clk),
	.d(\ex_csr_addr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_addr[1]~q ),
	.prn(vcc));
defparam \ex_csr_addr[1] .is_wysiwyg = "true";
defparam \ex_csr_addr[1] .power_up = "low";

cyclone10lp_lcell_comb \io_sw_r_ex_imm[1]~0 (
	.dataa(\ex_inst[16]~q ),
	.datab(\ex_csr_addr[1]~q ),
	.datac(gnd),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\io_sw_r_ex_imm[1]~0_combout ),
	.cout());
defparam \io_sw_r_ex_imm[1]~0 .lut_mask = 16'hAACC;
defparam \io_sw_r_ex_imm[1]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_op1~3 (
	.dataa(\ex_ctrl_alu_func~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal11~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_op1~3_combout ),
	.cout());
defparam \ex_ctrl_alu_op1~3 .lut_mask = 16'h00AA;
defparam \ex_ctrl_alu_op1~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_imm_type~15 (
	.dataa(\ex_ctrl_alu_op1~2_combout ),
	.datab(\ex_ctrl_mask_type~0_combout ),
	.datac(\Equal8~2_combout ),
	.datad(\ex_ctrl_alu_op1~3_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_imm_type~15_combout ),
	.cout());
defparam \ex_ctrl_imm_type~15 .lut_mask = 16'h0004;
defparam \ex_ctrl_imm_type~15 .sum_lutc_input = "datac";

dffeas \ex_ctrl_imm_type.010 (
	.clk(clk_clk),
	.d(\ex_ctrl_imm_type~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_imm_type.010~q ),
	.prn(vcc));
defparam \ex_ctrl_imm_type.010 .is_wysiwyg = "true";
defparam \ex_ctrl_imm_type.010 .power_up = "low";

cyclone10lp_lcell_comb \io_sw_r_ex_imm[1]~1 (
	.dataa(\ex_inst[8]~q ),
	.datab(\io_sw_r_ex_imm[1]~0_combout ),
	.datac(\ex_ctrl_imm_type.001~q ),
	.datad(\ex_ctrl_imm_type.010~q ),
	.cin(gnd),
	.combout(\io_sw_r_ex_imm[1]~1_combout ),
	.cout());
defparam \io_sw_r_ex_imm[1]~1 .lut_mask = 16'hAAAC;
defparam \io_sw_r_ex_imm[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_imm_type~16 (
	.dataa(\Equal5~0_combout ),
	.datab(\id_inst[4]~q ),
	.datac(gnd),
	.datad(\id_inst[6]~q ),
	.cin(gnd),
	.combout(\ex_ctrl_imm_type~16_combout ),
	.cout());
defparam \ex_ctrl_imm_type~16 .lut_mask = 16'h0088;
defparam \ex_ctrl_imm_type~16 .sum_lutc_input = "datac";

dffeas \ex_ctrl_imm_type.011 (
	.clk(clk_clk),
	.d(\ex_ctrl_imm_type~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\id_pc[7]~31_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_imm_type.011~q ),
	.prn(vcc));
defparam \ex_ctrl_imm_type.011 .is_wysiwyg = "true";
defparam \ex_ctrl_imm_type.011 .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~16 (
	.dataa(\io_sw_r_ex_imm[1]~1_combout ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\mem_imm~16_combout ),
	.cout());
defparam \mem_imm~16 .lut_mask = 16'h0088;
defparam \mem_imm~16 .sum_lutc_input = "datac";

dffeas \mem_imm[1] (
	.clk(clk_clk),
	.d(\mem_imm~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[1]~q ),
	.prn(vcc));
defparam \mem_imm[1] .is_wysiwyg = "true";
defparam \mem_imm[1] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[1]~2 (
	.dataa(gnd),
	.datab(\mem_imm[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\_T_3862[1]~2_combout ),
	.cout());
defparam \_T_3862[1]~2 .lut_mask = 16'hCCCC;
defparam \_T_3862[1]~2 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~5 (
	.dataa(\pc_cntr[0]~1_combout ),
	.datab(\csr|mepc[1]~q ),
	.datac(\pc_cntr[0]~0_combout ),
	.datad(mem_alu_out_1),
	.cin(gnd),
	.combout(\pc_cntr~5_combout ),
	.cout());
defparam \pc_cntr~5 .lut_mask = 16'hE5E0;
defparam \pc_cntr~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~6 (
	.dataa(\_T_3862[1]~2_combout ),
	.datab(\pc_cntr[0]~1_combout ),
	.datac(\pc_cntr~5_combout ),
	.datad(\csr|mtvec[1]~q ),
	.cin(gnd),
	.combout(\pc_cntr~6_combout ),
	.cout());
defparam \pc_cntr~6 .lut_mask = 16'hF838;
defparam \pc_cntr~6 .sum_lutc_input = "datac";

dffeas \pc_cntr[1] (
	.clk(clk_clk),
	.d(\pc_cntr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(\pc_cntr[0]~4_combout ),
	.q(\pc_cntr[1]~q ),
	.prn(vcc));
defparam \pc_cntr[1] .is_wysiwyg = "true";
defparam \pc_cntr[1] .power_up = "low";

cyclone10lp_lcell_comb \id_npc~1 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~1_combout ),
	.cout());
defparam \id_npc~1 .lut_mask = 16'h8080;
defparam \id_npc~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~4 (
	.dataa(id_pc_2),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~4_combout ),
	.cout());
defparam \ex_pc~4 .lut_mask = 16'h8080;
defparam \ex_pc~4 .sum_lutc_input = "datac";

dffeas \ex_pc[2] (
	.clk(clk_clk),
	.d(\ex_pc~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[2]~q ),
	.prn(vcc));
defparam \ex_pc[2] .is_wysiwyg = "true";
defparam \ex_pc[2] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~0 (
	.dataa(\ex_pc[2]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~0_combout ),
	.cout());
defparam \mem_pc~0 .lut_mask = 16'h8888;
defparam \mem_pc~0 .sum_lutc_input = "datac";

dffeas \mem_pc[2] (
	.clk(clk_clk),
	.d(\mem_pc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[2]~q ),
	.prn(vcc));
defparam \mem_pc[2] .is_wysiwyg = "true";
defparam \mem_pc[2] .power_up = "low";

cyclone10lp_lcell_comb \ex_inst~7 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~7_combout ),
	.cout());
defparam \ex_inst~7 .lut_mask = 16'h8080;
defparam \ex_inst~7 .sum_lutc_input = "datac";

dffeas \ex_inst[9] (
	.clk(clk_clk),
	.d(\ex_inst~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[9]~q ),
	.prn(vcc));
defparam \ex_inst[9] .is_wysiwyg = "true";
defparam \ex_inst[9] .power_up = "low";

cyclone10lp_lcell_comb \ex_inst~2 (
	.dataa(\id_inst[17]~q ),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~2_combout ),
	.cout());
defparam \ex_inst~2 .lut_mask = 16'h8080;
defparam \ex_inst~2 .sum_lutc_input = "datac";

dffeas \ex_inst[17] (
	.clk(clk_clk),
	.d(\ex_inst~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[17]~q ),
	.prn(vcc));
defparam \ex_inst[17] .is_wysiwyg = "true";
defparam \ex_inst[17] .power_up = "low";

cyclone10lp_lcell_comb \ex_csr_addr~2 (
	.dataa(\id_inst[22]~q ),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_csr_addr~2_combout ),
	.cout());
defparam \ex_csr_addr~2 .lut_mask = 16'h8080;
defparam \ex_csr_addr~2 .sum_lutc_input = "datac";

dffeas \ex_csr_addr[2] (
	.clk(clk_clk),
	.d(\ex_csr_addr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_addr[2]~q ),
	.prn(vcc));
defparam \ex_csr_addr[2] .is_wysiwyg = "true";
defparam \ex_csr_addr[2] .power_up = "low";

cyclone10lp_lcell_comb \io_sw_r_ex_imm[2]~5 (
	.dataa(\ex_inst[17]~q ),
	.datab(\ex_csr_addr[2]~q ),
	.datac(gnd),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\io_sw_r_ex_imm[2]~5_combout ),
	.cout());
defparam \io_sw_r_ex_imm[2]~5 .lut_mask = 16'hAACC;
defparam \io_sw_r_ex_imm[2]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_sw_r_ex_imm[2]~6 (
	.dataa(\ex_inst[9]~q ),
	.datab(\io_sw_r_ex_imm[2]~5_combout ),
	.datac(\ex_ctrl_imm_type.001~q ),
	.datad(\ex_ctrl_imm_type.010~q ),
	.cin(gnd),
	.combout(\io_sw_r_ex_imm[2]~6_combout ),
	.cout());
defparam \io_sw_r_ex_imm[2]~6 .lut_mask = 16'hAAAC;
defparam \io_sw_r_ex_imm[2]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~17 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\io_sw_r_ex_imm[2]~6_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\mem_imm~17_combout ),
	.cout());
defparam \mem_imm~17 .lut_mask = 16'h0088;
defparam \mem_imm~17 .sum_lutc_input = "datac";

dffeas \mem_imm[2] (
	.clk(clk_clk),
	.d(\mem_imm~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[2]~q ),
	.prn(vcc));
defparam \mem_imm[2] .is_wysiwyg = "true";
defparam \mem_imm[2] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[2]~4 (
	.dataa(\mem_pc[2]~q ),
	.datab(\mem_imm[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\_T_3862[2]~4_combout ),
	.cout(\_T_3862[2]~5 ));
defparam \_T_3862[2]~4 .lut_mask = 16'h6688;
defparam \_T_3862[2]~4 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr[19]~7 (
	.dataa(\Equal2~0_combout ),
	.datab(\mem_alu_cmp_out~q ),
	.datac(\mem_ctrl_br_type[0]~q ),
	.datad(\mem_ctrl_br_type[1]~q ),
	.cin(gnd),
	.combout(\pc_cntr[19]~7_combout ),
	.cout());
defparam \pc_cntr[19]~7 .lut_mask = 16'h1BBB;
defparam \pc_cntr[19]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr[19]~8 (
	.dataa(\mem_ctrl_br_type[0]~q ),
	.datab(\mem_ctrl_br_type[1]~q ),
	.datac(\mem_ctrl_br_type[2]~q ),
	.datad(\mem_ctrl_br_type[3]~q ),
	.cin(gnd),
	.combout(\pc_cntr[19]~8_combout ),
	.cout());
defparam \pc_cntr[19]~8 .lut_mask = 16'h000E;
defparam \pc_cntr[19]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \npc[2]~0 (
	.dataa(\pc_cntr[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\npc[2]~0_combout ),
	.cout(\npc[2]~1 ));
defparam \npc[2]~0 .lut_mask = 16'h55AA;
defparam \npc[2]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~9 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(mem_alu_out_2),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[2]~0_combout ),
	.cin(gnd),
	.combout(\pc_cntr~9_combout ),
	.cout());
defparam \pc_cntr~9 .lut_mask = 16'hDAD0;
defparam \pc_cntr~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~10 (
	.dataa(\_T_3862[2]~4_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~9_combout ),
	.datad(\csr|mepc[2]~q ),
	.cin(gnd),
	.combout(\pc_cntr~10_combout ),
	.cout());
defparam \pc_cntr~10 .lut_mask = 16'hF2C2;
defparam \pc_cntr~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~11 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~10_combout ),
	.datac(\csr|mtvec[2]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~11_combout ),
	.cout());
defparam \pc_cntr~11 .lut_mask = 16'h88A0;
defparam \pc_cntr~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr[19]~12 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(gnd),
	.datac(gnd),
	.datad(\csr|mcause[0]~6_combout ),
	.cin(gnd),
	.combout(\pc_cntr[19]~12_combout ),
	.cout());
defparam \pc_cntr[19]~12 .lut_mask = 16'hFF55;
defparam \pc_cntr[19]~12 .sum_lutc_input = "datac";

dffeas \pc_cntr[2] (
	.clk(clk_clk),
	.d(\pc_cntr~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[2]~q ),
	.prn(vcc));
defparam \pc_cntr[2] .is_wysiwyg = "true";
defparam \pc_cntr[2] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~1 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~1_combout ),
	.cout());
defparam \id_pc~1 .lut_mask = 16'h8080;
defparam \id_pc~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~5 (
	.dataa(id_pc_3),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~5_combout ),
	.cout());
defparam \ex_pc~5 .lut_mask = 16'h8080;
defparam \ex_pc~5 .sum_lutc_input = "datac";

dffeas \ex_pc[3] (
	.clk(clk_clk),
	.d(\ex_pc~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[3]~q ),
	.prn(vcc));
defparam \ex_pc[3] .is_wysiwyg = "true";
defparam \ex_pc[3] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~1 (
	.dataa(\ex_pc[3]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~1_combout ),
	.cout());
defparam \mem_pc~1 .lut_mask = 16'h8888;
defparam \mem_pc~1 .sum_lutc_input = "datac";

dffeas \mem_pc[3] (
	.clk(clk_clk),
	.d(\mem_pc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[3]~q ),
	.prn(vcc));
defparam \mem_pc[3] .is_wysiwyg = "true";
defparam \mem_pc[3] .power_up = "low";

cyclone10lp_lcell_comb \ex_inst~8 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[10]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~8_combout ),
	.cout());
defparam \ex_inst~8 .lut_mask = 16'h8080;
defparam \ex_inst~8 .sum_lutc_input = "datac";

dffeas \ex_inst[10] (
	.clk(clk_clk),
	.d(\ex_inst~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[10]~q ),
	.prn(vcc));
defparam \ex_inst[10] .is_wysiwyg = "true";
defparam \ex_inst[10] .power_up = "low";

cyclone10lp_lcell_comb \ex_inst~3 (
	.dataa(\id_inst[18]~q ),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~3_combout ),
	.cout());
defparam \ex_inst~3 .lut_mask = 16'h8080;
defparam \ex_inst~3 .sum_lutc_input = "datac";

dffeas \ex_inst[18] (
	.clk(clk_clk),
	.d(\ex_inst~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[18]~q ),
	.prn(vcc));
defparam \ex_inst[18] .is_wysiwyg = "true";
defparam \ex_inst[18] .power_up = "low";

cyclone10lp_lcell_comb \ex_csr_addr~3 (
	.dataa(\id_inst[23]~q ),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_csr_addr~3_combout ),
	.cout());
defparam \ex_csr_addr~3 .lut_mask = 16'h8080;
defparam \ex_csr_addr~3 .sum_lutc_input = "datac";

dffeas \ex_csr_addr[3] (
	.clk(clk_clk),
	.d(\ex_csr_addr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_addr[3]~q ),
	.prn(vcc));
defparam \ex_csr_addr[3] .is_wysiwyg = "true";
defparam \ex_csr_addr[3] .power_up = "low";

cyclone10lp_lcell_comb \io_sw_r_ex_imm[3]~7 (
	.dataa(\ex_inst[18]~q ),
	.datab(\ex_csr_addr[3]~q ),
	.datac(gnd),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\io_sw_r_ex_imm[3]~7_combout ),
	.cout());
defparam \io_sw_r_ex_imm[3]~7 .lut_mask = 16'hAACC;
defparam \io_sw_r_ex_imm[3]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_sw_r_ex_imm[3]~8 (
	.dataa(\ex_inst[10]~q ),
	.datab(\io_sw_r_ex_imm[3]~7_combout ),
	.datac(\ex_ctrl_imm_type.001~q ),
	.datad(\ex_ctrl_imm_type.010~q ),
	.cin(gnd),
	.combout(\io_sw_r_ex_imm[3]~8_combout ),
	.cout());
defparam \io_sw_r_ex_imm[3]~8 .lut_mask = 16'hAAAC;
defparam \io_sw_r_ex_imm[3]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~18 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\io_sw_r_ex_imm[3]~8_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\mem_imm~18_combout ),
	.cout());
defparam \mem_imm~18 .lut_mask = 16'h0088;
defparam \mem_imm~18 .sum_lutc_input = "datac";

dffeas \mem_imm[3] (
	.clk(clk_clk),
	.d(\mem_imm~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[3]~q ),
	.prn(vcc));
defparam \mem_imm[3] .is_wysiwyg = "true";
defparam \mem_imm[3] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[3]~6 (
	.dataa(\mem_pc[3]~q ),
	.datab(\mem_imm[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[2]~5 ),
	.combout(\_T_3862[3]~6_combout ),
	.cout(\_T_3862[3]~7 ));
defparam \_T_3862[3]~6 .lut_mask = 16'h9617;
defparam \_T_3862[3]~6 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \npc[3]~2 (
	.dataa(\pc_cntr[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[2]~1 ),
	.combout(\npc[3]~2_combout ),
	.cout(\npc[3]~3 ));
defparam \npc[3]~2 .lut_mask = 16'h5A5F;
defparam \npc[3]~2 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~13 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[3]~6_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[3]~2_combout ),
	.cin(gnd),
	.combout(\pc_cntr~13_combout ),
	.cout());
defparam \pc_cntr~13 .lut_mask = 16'h5E0E;
defparam \pc_cntr~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~14 (
	.dataa(mem_alu_out_3),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~13_combout ),
	.datad(\csr|mepc[3]~q ),
	.cin(gnd),
	.combout(\pc_cntr~14_combout ),
	.cout());
defparam \pc_cntr~14 .lut_mask = 16'hF838;
defparam \pc_cntr~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~15 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~14_combout ),
	.datac(\csr|mtvec[3]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~15_combout ),
	.cout());
defparam \pc_cntr~15 .lut_mask = 16'h88A0;
defparam \pc_cntr~15 .sum_lutc_input = "datac";

dffeas \pc_cntr[3] (
	.clk(clk_clk),
	.d(\pc_cntr~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[3]~q ),
	.prn(vcc));
defparam \pc_cntr[3] .is_wysiwyg = "true";
defparam \pc_cntr[3] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~2 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~2_combout ),
	.cout());
defparam \id_pc~2 .lut_mask = 16'h8080;
defparam \id_pc~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~0 (
	.dataa(id_pc_4),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~0_combout ),
	.cout());
defparam \ex_pc~0 .lut_mask = 16'h8080;
defparam \ex_pc~0 .sum_lutc_input = "datac";

dffeas \ex_pc[4] (
	.clk(clk_clk),
	.d(\ex_pc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[4]~q ),
	.prn(vcc));
defparam \ex_pc[4] .is_wysiwyg = "true";
defparam \ex_pc[4] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~2 (
	.dataa(\ex_pc[4]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~2_combout ),
	.cout());
defparam \mem_pc~2 .lut_mask = 16'h8888;
defparam \mem_pc~2 .sum_lutc_input = "datac";

dffeas \mem_pc[4] (
	.clk(clk_clk),
	.d(\mem_pc~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[4]~q ),
	.prn(vcc));
defparam \mem_pc[4] .is_wysiwyg = "true";
defparam \mem_pc[4] .power_up = "low";

cyclone10lp_lcell_comb \ex_inst~9 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[11]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~9_combout ),
	.cout());
defparam \ex_inst~9 .lut_mask = 16'h8080;
defparam \ex_inst~9 .sum_lutc_input = "datac";

dffeas \ex_inst[11] (
	.clk(clk_clk),
	.d(\ex_inst~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[11]~q ),
	.prn(vcc));
defparam \ex_inst[11] .is_wysiwyg = "true";
defparam \ex_inst[11] .power_up = "low";

cyclone10lp_lcell_comb \ex_inst~4 (
	.dataa(\id_inst[19]~q ),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~4_combout ),
	.cout());
defparam \ex_inst~4 .lut_mask = 16'h8080;
defparam \ex_inst~4 .sum_lutc_input = "datac";

dffeas \ex_inst[19] (
	.clk(clk_clk),
	.d(\ex_inst~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[19]~q ),
	.prn(vcc));
defparam \ex_inst[19] .is_wysiwyg = "true";
defparam \ex_inst[19] .power_up = "low";

cyclone10lp_lcell_comb \ex_csr_addr~4 (
	.dataa(\id_inst[24]~q ),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_csr_addr~4_combout ),
	.cout());
defparam \ex_csr_addr~4 .lut_mask = 16'h8080;
defparam \ex_csr_addr~4 .sum_lutc_input = "datac";

dffeas \ex_csr_addr[4] (
	.clk(clk_clk),
	.d(\ex_csr_addr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_addr[4]~q ),
	.prn(vcc));
defparam \ex_csr_addr[4] .is_wysiwyg = "true";
defparam \ex_csr_addr[4] .power_up = "low";

cyclone10lp_lcell_comb \io_sw_r_ex_imm[4]~3 (
	.dataa(\ex_inst[19]~q ),
	.datab(\ex_csr_addr[4]~q ),
	.datac(gnd),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\io_sw_r_ex_imm[4]~3_combout ),
	.cout());
defparam \io_sw_r_ex_imm[4]~3 .lut_mask = 16'hAACC;
defparam \io_sw_r_ex_imm[4]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_sw_r_ex_imm[4]~4 (
	.dataa(\ex_inst[11]~q ),
	.datab(\io_sw_r_ex_imm[4]~3_combout ),
	.datac(\ex_ctrl_imm_type.001~q ),
	.datad(\ex_ctrl_imm_type.010~q ),
	.cin(gnd),
	.combout(\io_sw_r_ex_imm[4]~4_combout ),
	.cout());
defparam \io_sw_r_ex_imm[4]~4 .lut_mask = 16'hAAAC;
defparam \io_sw_r_ex_imm[4]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~19 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\io_sw_r_ex_imm[4]~4_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\mem_imm~19_combout ),
	.cout());
defparam \mem_imm~19 .lut_mask = 16'h0088;
defparam \mem_imm~19 .sum_lutc_input = "datac";

dffeas \mem_imm[4] (
	.clk(clk_clk),
	.d(\mem_imm~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[4]~q ),
	.prn(vcc));
defparam \mem_imm[4] .is_wysiwyg = "true";
defparam \mem_imm[4] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[4]~8 (
	.dataa(\mem_pc[4]~q ),
	.datab(\mem_imm[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[3]~7 ),
	.combout(\_T_3862[4]~8_combout ),
	.cout(\_T_3862[4]~9 ));
defparam \_T_3862[4]~8 .lut_mask = 16'h698E;
defparam \_T_3862[4]~8 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \ex_ctrl_alu_op2~6 (
	.dataa(\ex_ctrl_alu_op2~5_combout ),
	.datab(\ex_ctrl_mask_type~0_combout ),
	.datac(\_T_3083~0_combout ),
	.datad(\ex_ctrl_csr_cmd~9_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_op2~6_combout ),
	.cout());
defparam \ex_ctrl_alu_op2~6 .lut_mask = 16'h8000;
defparam \ex_ctrl_alu_op2~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_op2~7 (
	.dataa(\ex_ctrl_imm_type~15_combout ),
	.datab(gnd),
	.datac(\ex_ctrl_alu_op2~6_combout ),
	.datad(\ex_ctrl_csr_cmd~10_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_op2~7_combout ),
	.cout());
defparam \ex_ctrl_alu_op2~7 .lut_mask = 16'h0AFA;
defparam \ex_ctrl_alu_op2~7 .sum_lutc_input = "datac";

dffeas \ex_ctrl_alu_op2.01 (
	.clk(clk_clk),
	.d(\ex_ctrl_alu_op2~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_alu_op2.01~q ),
	.prn(vcc));
defparam \ex_ctrl_alu_op2.01 .is_wysiwyg = "true";
defparam \ex_ctrl_alu_op2.01 .power_up = "low";

cyclone10lp_lcell_comb \ex_ctrl_alu_op2~8 (
	.dataa(gnd),
	.datab(\ex_ctrl_alu_op2~6_combout ),
	.datac(\ex_ctrl_imm_type~15_combout ),
	.datad(\ex_ctrl_imm_type~13_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_op2~8_combout ),
	.cout());
defparam \ex_ctrl_alu_op2~8 .lut_mask = 16'hFC30;
defparam \ex_ctrl_alu_op2~8 .sum_lutc_input = "datac";

dffeas \ex_ctrl_alu_op2.10 (
	.clk(clk_clk),
	.d(\ex_ctrl_alu_op2~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_alu_op2.10~q ),
	.prn(vcc));
defparam \ex_ctrl_alu_op2.10 .is_wysiwyg = "true";
defparam \ex_ctrl_alu_op2.10 .power_up = "low";

cyclone10lp_lcell_comb \csr_io_alu_op2[1]~0 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(gnd),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\csr_io_alu_op2[1]~0_combout ),
	.cout());
defparam \csr_io_alu_op2[1]~0 .lut_mask = 16'h88BB;
defparam \csr_io_alu_op2[1]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_csr_cmd~4 (
	.dataa(gnd),
	.datab(\id_inst[4]~q ),
	.datac(\id_inst[6]~q ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\ex_csr_cmd~4_combout ),
	.cout());
defparam \ex_csr_cmd~4 .lut_mask = 16'h3FFF;
defparam \ex_csr_cmd~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~5 (
	.dataa(\id_inst[25]~q ),
	.datab(gnd),
	.datac(\id_inst[14]~q ),
	.datad(\Equal29~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~5_combout ),
	.cout());
defparam \ex_ctrl_alu_func~5 .lut_mask = 16'h0AFF;
defparam \ex_ctrl_alu_func~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_csr_cmd~11 (
	.dataa(\ex_ctrl_alu_func~5_combout ),
	.datab(\_T_3083~0_combout ),
	.datac(\ex_ctrl_csr_cmd~10_combout ),
	.datad(\Equal31~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_csr_cmd~11_combout ),
	.cout());
defparam \ex_ctrl_csr_cmd~11 .lut_mask = 16'h0080;
defparam \ex_ctrl_csr_cmd~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal45~0 (
	.dataa(\id_inst[4]~q ),
	.datab(\id_inst[6]~q ),
	.datac(\Equal10~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal45~0_combout ),
	.cout());
defparam \Equal45~0 .lut_mask = 16'h8080;
defparam \Equal45~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_csr_cmd~12 (
	.dataa(\ex_ctrl_csr_cmd~9_combout ),
	.datab(\ex_ctrl_imm_type~13_combout ),
	.datac(\ex_ctrl_csr_cmd~11_combout ),
	.datad(\Equal45~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_csr_cmd~12_combout ),
	.cout());
defparam \ex_ctrl_csr_cmd~12 .lut_mask = 16'h0080;
defparam \ex_ctrl_csr_cmd~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal48~4 (
	.dataa(\Equal8~0_combout ),
	.datab(\Equal48~3_combout ),
	.datac(\Equal29~0_combout ),
	.datad(\id_inst[21]~q ),
	.cin(gnd),
	.combout(\Equal48~4_combout ),
	.cout());
defparam \Equal48~4 .lut_mask = 16'h0080;
defparam \Equal48~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_wb_sel~10 (
	.dataa(\id_inst[20]~q ),
	.datab(gnd),
	.datac(\Equal48~4_combout ),
	.datad(\Equal49~3_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_wb_sel~10_combout ),
	.cout());
defparam \ex_ctrl_wb_sel~10 .lut_mask = 16'h00AF;
defparam \ex_ctrl_wb_sel~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal50~0 (
	.dataa(\Equal49~2_combout ),
	.datab(gnd),
	.datac(\id_inst[21]~q ),
	.datad(\id_inst[29]~q ),
	.cin(gnd),
	.combout(\Equal50~0_combout ),
	.cout());
defparam \Equal50~0 .lut_mask = 16'h000A;
defparam \Equal50~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_csr_cmd~13 (
	.dataa(\ex_csr_cmd~4_combout ),
	.datab(\ex_ctrl_csr_cmd~12_combout ),
	.datac(\ex_ctrl_wb_sel~10_combout ),
	.datad(\Equal50~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_csr_cmd~13_combout ),
	.cout());
defparam \ex_ctrl_csr_cmd~13 .lut_mask = 16'h0080;
defparam \ex_ctrl_csr_cmd~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal51~0 (
	.dataa(\id_inst[20]~q ),
	.datab(\Equal48~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal51~0_combout ),
	.cout());
defparam \Equal51~0 .lut_mask = 16'h8888;
defparam \Equal51~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_csr_cmd~16 (
	.dataa(\ex_ctrl_csr_cmd~14_combout ),
	.datab(\ex_ctrl_csr_cmd~13_combout ),
	.datac(\Equal51~0_combout ),
	.datad(\ex_ctrl_mask_type~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_csr_cmd~16_combout ),
	.cout());
defparam \ex_ctrl_csr_cmd~16 .lut_mask = 16'hD100;
defparam \ex_ctrl_csr_cmd~16 .sum_lutc_input = "datac";

dffeas \ex_ctrl_csr_cmd.000 (
	.clk(clk_clk),
	.d(\ex_ctrl_csr_cmd~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_csr_cmd.000~q ),
	.prn(vcc));
defparam \ex_ctrl_csr_cmd.000 .is_wysiwyg = "true";
defparam \ex_ctrl_csr_cmd.000 .power_up = "low";

cyclone10lp_lcell_comb \mem_ctrl_csr_cmd~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\mem_ctrl_mem_wr~7_combout ),
	.datad(\ex_ctrl_csr_cmd.000~q ),
	.cin(gnd),
	.combout(\mem_ctrl_csr_cmd~14_combout ),
	.cout());
defparam \mem_ctrl_csr_cmd~14 .lut_mask = 16'hF000;
defparam \mem_ctrl_csr_cmd~14 .sum_lutc_input = "datac";

dffeas \mem_ctrl_csr_cmd.000 (
	.clk(clk_clk),
	.d(\mem_ctrl_csr_cmd~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_ctrl_csr_cmd.000~q ),
	.prn(vcc));
defparam \mem_ctrl_csr_cmd.000 .is_wysiwyg = "true";
defparam \mem_ctrl_csr_cmd.000 .power_up = "low";

cyclone10lp_lcell_comb \mem_reg_waddr~1 (
	.dataa(\ex_inst[8]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_reg_waddr~1_combout ),
	.cout());
defparam \mem_reg_waddr~1 .lut_mask = 16'h8888;
defparam \mem_reg_waddr~1 .sum_lutc_input = "datac";

dffeas \mem_reg_waddr[1] (
	.clk(clk_clk),
	.d(\mem_reg_waddr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_reg_waddr[1]~q ),
	.prn(vcc));
defparam \mem_reg_waddr[1] .is_wysiwyg = "true";
defparam \mem_reg_waddr[1] .power_up = "low";

cyclone10lp_lcell_comb \mem_reg_waddr~0 (
	.dataa(\ex_inst[7]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_reg_waddr~0_combout ),
	.cout());
defparam \mem_reg_waddr~0 .lut_mask = 16'h8888;
defparam \mem_reg_waddr~0 .sum_lutc_input = "datac";

dffeas \mem_reg_waddr[0] (
	.clk(clk_clk),
	.d(\mem_reg_waddr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_reg_waddr[0]~q ),
	.prn(vcc));
defparam \mem_reg_waddr[0] .is_wysiwyg = "true";
defparam \mem_reg_waddr[0] .power_up = "low";

cyclone10lp_lcell_comb \_T_3681~0 (
	.dataa(\ex_csr_addr[0]~q ),
	.datab(\ex_csr_addr[1]~q ),
	.datac(\mem_reg_waddr[1]~q ),
	.datad(\mem_reg_waddr[0]~q ),
	.cin(gnd),
	.combout(\_T_3681~0_combout ),
	.cout());
defparam \_T_3681~0 .lut_mask = 16'h8241;
defparam \_T_3681~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_reg_waddr~3 (
	.dataa(\ex_inst[10]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_reg_waddr~3_combout ),
	.cout());
defparam \mem_reg_waddr~3 .lut_mask = 16'h8888;
defparam \mem_reg_waddr~3 .sum_lutc_input = "datac";

dffeas \mem_reg_waddr[3] (
	.clk(clk_clk),
	.d(\mem_reg_waddr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_reg_waddr[3]~q ),
	.prn(vcc));
defparam \mem_reg_waddr[3] .is_wysiwyg = "true";
defparam \mem_reg_waddr[3] .power_up = "low";

cyclone10lp_lcell_comb \mem_reg_waddr~2 (
	.dataa(\ex_inst[9]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_reg_waddr~2_combout ),
	.cout());
defparam \mem_reg_waddr~2 .lut_mask = 16'h8888;
defparam \mem_reg_waddr~2 .sum_lutc_input = "datac";

dffeas \mem_reg_waddr[2] (
	.clk(clk_clk),
	.d(\mem_reg_waddr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_reg_waddr[2]~q ),
	.prn(vcc));
defparam \mem_reg_waddr[2] .is_wysiwyg = "true";
defparam \mem_reg_waddr[2] .power_up = "low";

cyclone10lp_lcell_comb \_T_3681~1 (
	.dataa(\ex_csr_addr[2]~q ),
	.datab(\ex_csr_addr[3]~q ),
	.datac(\mem_reg_waddr[3]~q ),
	.datad(\mem_reg_waddr[2]~q ),
	.cin(gnd),
	.combout(\_T_3681~1_combout ),
	.cout());
defparam \_T_3681~1 .lut_mask = 16'h8241;
defparam \_T_3681~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3681~2 (
	.dataa(\_T_3681~0_combout ),
	.datab(\_T_3681~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\_T_3681~2_combout ),
	.cout());
defparam \_T_3681~2 .lut_mask = 16'h8888;
defparam \_T_3681~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_reg_waddr~4 (
	.dataa(\ex_inst[11]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_reg_waddr~4_combout ),
	.cout());
defparam \mem_reg_waddr~4 .lut_mask = 16'h8888;
defparam \mem_reg_waddr~4 .sum_lutc_input = "datac";

dffeas \mem_reg_waddr[4] (
	.clk(clk_clk),
	.d(\mem_reg_waddr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_reg_waddr[4]~q ),
	.prn(vcc));
defparam \mem_reg_waddr[4] .is_wysiwyg = "true";
defparam \mem_reg_waddr[4] .power_up = "low";

cyclone10lp_lcell_comb \Equal63~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\mem_reg_waddr[4]~q ),
	.datad(\ex_csr_addr[4]~q ),
	.cin(gnd),
	.combout(\Equal63~0_combout ),
	.cout());
defparam \Equal63~0 .lut_mask = 16'h0FF0;
defparam \Equal63~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\ex_csr_addr[0]~q ),
	.datad(\ex_csr_addr[1]~q ),
	.cin(gnd),
	.combout(\Equal62~0_combout ),
	.cout());
defparam \Equal62~0 .lut_mask = 16'h000F;
defparam \Equal62~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal62~1 (
	.dataa(\Equal62~0_combout ),
	.datab(\ex_csr_addr[4]~q ),
	.datac(\ex_csr_addr[2]~q ),
	.datad(\ex_csr_addr[3]~q ),
	.cin(gnd),
	.combout(\Equal62~1_combout ),
	.cout());
defparam \Equal62~1 .lut_mask = 16'h0002;
defparam \Equal62~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3681~3 (
	.dataa(\mem_ctrl_csr_cmd.000~q ),
	.datab(\_T_3681~2_combout ),
	.datac(\Equal63~0_combout ),
	.datad(\Equal62~1_combout ),
	.cin(gnd),
	.combout(\_T_3681~3_combout ),
	.cout());
defparam \_T_3681~3 .lut_mask = 16'h0008;
defparam \_T_3681~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_csr_data~25 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[4]~142_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~25_combout ),
	.cout());
defparam \mem_csr_data~25 .lut_mask = 16'h8888;
defparam \mem_csr_data~25 .sum_lutc_input = "datac";

dffeas \mem_csr_data[4] (
	.clk(clk_clk),
	.d(\mem_csr_data~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[4]~q ),
	.prn(vcc));
defparam \mem_csr_data[4] .is_wysiwyg = "true";
defparam \mem_csr_data[4] .power_up = "low";

cyclone10lp_lcell_comb \ex_ctrl_rf_wen~0 (
	.dataa(\Equal5~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\ex_ctrl_rf_wen~0_combout ),
	.cout());
defparam \ex_ctrl_rf_wen~0 .lut_mask = 16'hAAFF;
defparam \ex_ctrl_rf_wen~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_op1~4 (
	.dataa(\ex_ctrl_alu_func~33_combout ),
	.datab(\ex_csr_cmd~4_combout ),
	.datac(gnd),
	.datad(\Equal8~2_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_op1~4_combout ),
	.cout());
defparam \ex_ctrl_alu_op1~4 .lut_mask = 16'h0088;
defparam \ex_ctrl_alu_op1~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_op1~5 (
	.dataa(\_T_1778~combout ),
	.datab(\ex_ctrl_csr_cmd~11_combout ),
	.datac(\ex_ctrl_alu_op1~4_combout ),
	.datad(\Equal45~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_op1~5_combout ),
	.cout());
defparam \ex_ctrl_alu_op1~5 .lut_mask = 16'h0080;
defparam \ex_ctrl_alu_op1~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_rf_wen~1 (
	.dataa(\ex_ctrl_rf_wen~0_combout ),
	.datab(\ex_ctrl_alu_op1~2_combout ),
	.datac(\ex_ctrl_imm_type~13_combout ),
	.datad(\ex_ctrl_alu_op1~5_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_rf_wen~1_combout ),
	.cout());
defparam \ex_ctrl_rf_wen~1 .lut_mask = 16'hEFFF;
defparam \ex_ctrl_rf_wen~1 .sum_lutc_input = "datac";

dffeas ex_ctrl_rf_wen(
	.clk(clk_clk),
	.d(\ex_ctrl_rf_wen~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_rf_wen~q ),
	.prn(vcc));
defparam ex_ctrl_rf_wen.is_wysiwyg = "true";
defparam ex_ctrl_rf_wen.power_up = "low";

cyclone10lp_lcell_comb \mem_ctrl_rf_wen~0 (
	.dataa(\ex_ctrl_rf_wen~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_ctrl_rf_wen~0_combout ),
	.cout());
defparam \mem_ctrl_rf_wen~0 .lut_mask = 16'hAAFF;
defparam \mem_ctrl_rf_wen~0 .sum_lutc_input = "datac";

dffeas mem_ctrl_rf_wen(
	.clk(clk_clk),
	.d(\mem_ctrl_rf_wen~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_ctrl_rf_wen~q ),
	.prn(vcc));
defparam mem_ctrl_rf_wen.is_wysiwyg = "true";
defparam mem_ctrl_rf_wen.power_up = "low";

cyclone10lp_lcell_comb \_T_3686~0 (
	.dataa(\_T_3681~2_combout ),
	.datab(\mem_ctrl_rf_wen~q ),
	.datac(\Equal63~0_combout ),
	.datad(\Equal62~1_combout ),
	.cin(gnd),
	.combout(\_T_3686~0_combout ),
	.cout());
defparam \_T_3686~0 .lut_mask = 16'h0008;
defparam \_T_3686~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_rs_1[23]~0 (
	.dataa(\id_inst[20]~q ),
	.datab(\id_inst[24]~q ),
	.datac(\id_inst[22]~q ),
	.datad(\id_inst[23]~q ),
	.cin(gnd),
	.combout(\ex_rs_1[23]~0_combout ),
	.cout());
defparam \ex_rs_1[23]~0 .lut_mask = 16'hFFFE;
defparam \ex_rs_1[23]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_rs_1[23]~1 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[21]~q ),
	.datad(\ex_rs_1[23]~0_combout ),
	.cin(gnd),
	.combout(\ex_rs_1[23]~1_combout ),
	.cout());
defparam \ex_rs_1[23]~1 .lut_mask = 16'h8880;
defparam \ex_rs_1[23]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_ctrl_rf_wen~0 (
	.dataa(\mem_ctrl_rf_wen~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\wb_ctrl_rf_wen~0_combout ),
	.cout());
defparam \wb_ctrl_rf_wen~0 .lut_mask = 16'hAAFF;
defparam \wb_ctrl_rf_wen~0 .sum_lutc_input = "datac";

dffeas wb_ctrl_rf_wen(
	.clk(clk_clk),
	.d(\wb_ctrl_rf_wen~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_ctrl_rf_wen~q ),
	.prn(vcc));
defparam wb_ctrl_rf_wen.is_wysiwyg = "true";
defparam wb_ctrl_rf_wen.power_up = "low";

cyclone10lp_lcell_comb \wb_reg_waddr~4 (
	.dataa(\mem_reg_waddr[4]~q ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_reg_waddr~4_combout ),
	.cout());
defparam \wb_reg_waddr~4 .lut_mask = 16'h8888;
defparam \wb_reg_waddr~4 .sum_lutc_input = "datac";

dffeas \wb_reg_waddr[4] (
	.clk(clk_clk),
	.d(\wb_reg_waddr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_reg_waddr[4]~q ),
	.prn(vcc));
defparam \wb_reg_waddr[4] .is_wysiwyg = "true";
defparam \wb_reg_waddr[4] .power_up = "low";

cyclone10lp_lcell_comb \wb_reg_waddr~0 (
	.dataa(\mem_reg_waddr[0]~q ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_reg_waddr~0_combout ),
	.cout());
defparam \wb_reg_waddr~0 .lut_mask = 16'h8888;
defparam \wb_reg_waddr~0 .sum_lutc_input = "datac";

dffeas \wb_reg_waddr[0] (
	.clk(clk_clk),
	.d(\wb_reg_waddr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_reg_waddr[0]~q ),
	.prn(vcc));
defparam \wb_reg_waddr[0] .is_wysiwyg = "true";
defparam \wb_reg_waddr[0] .power_up = "low";

cyclone10lp_lcell_comb \wb_reg_waddr~1 (
	.dataa(\mem_reg_waddr[1]~q ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_reg_waddr~1_combout ),
	.cout());
defparam \wb_reg_waddr~1 .lut_mask = 16'h8888;
defparam \wb_reg_waddr~1 .sum_lutc_input = "datac";

dffeas \wb_reg_waddr[1] (
	.clk(clk_clk),
	.d(\wb_reg_waddr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_reg_waddr[1]~q ),
	.prn(vcc));
defparam \wb_reg_waddr[1] .is_wysiwyg = "true";
defparam \wb_reg_waddr[1] .power_up = "low";

cyclone10lp_lcell_comb \wb_reg_waddr~2 (
	.dataa(\mem_reg_waddr[2]~q ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_reg_waddr~2_combout ),
	.cout());
defparam \wb_reg_waddr~2 .lut_mask = 16'h8888;
defparam \wb_reg_waddr~2 .sum_lutc_input = "datac";

dffeas \wb_reg_waddr[2] (
	.clk(clk_clk),
	.d(\wb_reg_waddr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_reg_waddr[2]~q ),
	.prn(vcc));
defparam \wb_reg_waddr[2] .is_wysiwyg = "true";
defparam \wb_reg_waddr[2] .power_up = "low";

cyclone10lp_lcell_comb \wb_reg_waddr~3 (
	.dataa(\mem_reg_waddr[3]~q ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_reg_waddr~3_combout ),
	.cout());
defparam \wb_reg_waddr~3 .lut_mask = 16'h8888;
defparam \wb_reg_waddr~3 .sum_lutc_input = "datac";

dffeas \wb_reg_waddr[3] (
	.clk(clk_clk),
	.d(\wb_reg_waddr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_reg_waddr[3]~q ),
	.prn(vcc));
defparam \wb_reg_waddr[3] .is_wysiwyg = "true";
defparam \wb_reg_waddr[3] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_en~0 (
	.dataa(\wb_reg_waddr[0]~q ),
	.datab(\wb_reg_waddr[1]~q ),
	.datac(\wb_reg_waddr[2]~q ),
	.datad(\wb_reg_waddr[3]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_en~0_combout ),
	.cout());
defparam \_T_3543__T_3854_en~0 .lut_mask = 16'hFFFE;
defparam \_T_3543__T_3854_en~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3543__T_3854_en~1 (
	.dataa(\wb_ctrl_rf_wen~q ),
	.datab(\wb_reg_waddr[4]~q ),
	.datac(\_T_3543__T_3854_en~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\_T_3543__T_3854_en~1_combout ),
	.cout());
defparam \_T_3543__T_3854_en~1 .lut_mask = 16'hA8A8;
defparam \_T_3543__T_3854_en~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_csr_data~18 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~18_combout ),
	.cout());
defparam \wb_csr_data~18 .lut_mask = 16'h8888;
defparam \wb_csr_data~18 .sum_lutc_input = "datac";

dffeas \wb_csr_data[4] (
	.clk(clk_clk),
	.d(\wb_csr_data~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[4]~q ),
	.prn(vcc));
defparam \wb_csr_data[4] .is_wysiwyg = "true";
defparam \wb_csr_data[4] .power_up = "low";

cyclone10lp_lcell_comb \wb_ctrl_wb_sel~14 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(mem_ctrl_mem_wr01),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_ctrl_wb_sel~14_combout ),
	.cout());
defparam \wb_ctrl_wb_sel~14 .lut_mask = 16'h8888;
defparam \wb_ctrl_wb_sel~14 .sum_lutc_input = "datac";

dffeas \wb_ctrl_wb_sel.10 (
	.clk(clk_clk),
	.d(\wb_ctrl_wb_sel~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_ctrl_wb_sel.10~q ),
	.prn(vcc));
defparam \wb_ctrl_wb_sel.10 .is_wysiwyg = "true";
defparam \wb_ctrl_wb_sel.10 .power_up = "low";

cyclone10lp_lcell_comb \ex_ctrl_wb_sel~11 (
	.dataa(\ex_ctrl_imm_type~13_combout ),
	.datab(\ex_csr_cmd~4_combout ),
	.datac(gnd),
	.datad(\Equal45~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_wb_sel~11_combout ),
	.cout());
defparam \ex_ctrl_wb_sel~11 .lut_mask = 16'h0088;
defparam \ex_ctrl_wb_sel~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_wb_sel~18 (
	.dataa(\ex_ctrl_wb_sel~10_combout ),
	.datab(\Equal50~0_combout ),
	.datac(\ex_ctrl_wb_sel~11_combout ),
	.datad(\ex_ctrl_csr_cmd~14_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_wb_sel~18_combout ),
	.cout());
defparam \ex_ctrl_wb_sel~18 .lut_mask = 16'h008F;
defparam \ex_ctrl_wb_sel~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_wb_sel~19 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\ex_ctrl_wb_sel~18_combout ),
	.datad(\Equal5~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_wb_sel~19_combout ),
	.cout());
defparam \ex_ctrl_wb_sel~19 .lut_mask = 16'h0080;
defparam \ex_ctrl_wb_sel~19 .sum_lutc_input = "datac";

dffeas \ex_ctrl_wb_sel.11 (
	.clk(clk_clk),
	.d(\ex_ctrl_wb_sel~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_wb_sel.11~q ),
	.prn(vcc));
defparam \ex_ctrl_wb_sel.11 .is_wysiwyg = "true";
defparam \ex_ctrl_wb_sel.11 .power_up = "low";

cyclone10lp_lcell_comb \mem_ctrl_wb_sel~13 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_ctrl_wb_sel.11~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_ctrl_wb_sel~13_combout ),
	.cout());
defparam \mem_ctrl_wb_sel~13 .lut_mask = 16'h8888;
defparam \mem_ctrl_wb_sel~13 .sum_lutc_input = "datac";

dffeas \mem_ctrl_wb_sel.11 (
	.clk(clk_clk),
	.d(\mem_ctrl_wb_sel~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_ctrl_wb_sel.11~q ),
	.prn(vcc));
defparam \mem_ctrl_wb_sel.11 .is_wysiwyg = "true";
defparam \mem_ctrl_wb_sel.11 .power_up = "low";

cyclone10lp_lcell_comb \wb_ctrl_wb_sel~13 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_ctrl_wb_sel.11~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_ctrl_wb_sel~13_combout ),
	.cout());
defparam \wb_ctrl_wb_sel~13 .lut_mask = 16'h8888;
defparam \wb_ctrl_wb_sel~13 .sum_lutc_input = "datac";

dffeas \wb_ctrl_wb_sel.11 (
	.clk(clk_clk),
	.d(\wb_ctrl_wb_sel~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_ctrl_wb_sel.11~q ),
	.prn(vcc));
defparam \wb_ctrl_wb_sel.11 .is_wysiwyg = "true";
defparam \wb_ctrl_wb_sel.11 .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[23]~2 (
	.dataa(\wb_ctrl_wb_sel.10~q ),
	.datab(\wb_ctrl_wb_sel.11~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[23]~2_combout ),
	.cout());
defparam \_T_3543__T_3854_data[23]~2 .lut_mask = 16'hEEEE;
defparam \_T_3543__T_3854_data[23]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \npc[4]~4 (
	.dataa(\pc_cntr[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[3]~3 ),
	.combout(\npc[4]~4_combout ),
	.cout(\npc[4]~5 ));
defparam \npc[4]~4 .lut_mask = 16'hA50A;
defparam \npc[4]~4 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~18 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[4]~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~18_combout ),
	.cout());
defparam \id_npc~18 .lut_mask = 16'h8080;
defparam \id_npc~18 .sum_lutc_input = "datac";

dffeas \id_npc[4] (
	.clk(clk_clk),
	.d(\id_npc~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[4]~q ),
	.prn(vcc));
defparam \id_npc[4] .is_wysiwyg = "true";
defparam \id_npc[4] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~18 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~18_combout ),
	.cout());
defparam \ex_npc~18 .lut_mask = 16'h8080;
defparam \ex_npc~18 .sum_lutc_input = "datac";

dffeas \ex_npc[4] (
	.clk(clk_clk),
	.d(\ex_npc~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[4]~q ),
	.prn(vcc));
defparam \ex_npc[4] .is_wysiwyg = "true";
defparam \ex_npc[4] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~16 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~16_combout ),
	.cout());
defparam \mem_npc~16 .lut_mask = 16'h8888;
defparam \mem_npc~16 .sum_lutc_input = "datac";

dffeas \mem_npc[4] (
	.clk(clk_clk),
	.d(\mem_npc~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[4]~q ),
	.prn(vcc));
defparam \mem_npc[4] .is_wysiwyg = "true";
defparam \mem_npc[4] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~16 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~16_combout ),
	.cout());
defparam \wb_npc~16 .lut_mask = 16'h8888;
defparam \wb_npc~16 .sum_lutc_input = "datac";

dffeas \wb_npc[4] (
	.clk(clk_clk),
	.d(\wb_npc~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[4]~q ),
	.prn(vcc));
defparam \wb_npc[4] .is_wysiwyg = "true";
defparam \wb_npc[4] .power_up = "low";

cyclone10lp_lcell_comb \ex_ctrl_wb_sel~13 (
	.dataa(\ex_ctrl_alu_func~33_combout ),
	.datab(\ex_ctrl_csr_cmd~11_combout ),
	.datac(\ex_ctrl_wb_sel~11_combout ),
	.datad(\ex_ctrl_imm_type~12_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_wb_sel~13_combout ),
	.cout());
defparam \ex_ctrl_wb_sel~13 .lut_mask = 16'h80AA;
defparam \ex_ctrl_wb_sel~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_wb_sel~14 (
	.dataa(\Equal8~2_combout ),
	.datab(\Equal7~0_combout ),
	.datac(\Equal53~0_combout ),
	.datad(\id_inst[4]~q ),
	.cin(gnd),
	.combout(\ex_ctrl_wb_sel~14_combout ),
	.cout());
defparam \ex_ctrl_wb_sel~14 .lut_mask = 16'hAAEA;
defparam \ex_ctrl_wb_sel~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_wb_sel~15 (
	.dataa(\ex_ctrl_wb_sel~13_combout ),
	.datab(\ex_ctrl_wb_sel~14_combout ),
	.datac(\ex_ctrl_alu_op1~3_combout ),
	.datad(\Equal6~3_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_wb_sel~15_combout ),
	.cout());
defparam \ex_ctrl_wb_sel~15 .lut_mask = 16'h00EF;
defparam \ex_ctrl_wb_sel~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_wb_sel~12 (
	.dataa(\ex_ctrl_csr_cmd~9_combout ),
	.datab(\ex_ctrl_csr_cmd~11_combout ),
	.datac(\ex_ctrl_wb_sel~11_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_ctrl_wb_sel~12_combout ),
	.cout());
defparam \ex_ctrl_wb_sel~12 .lut_mask = 16'h8080;
defparam \ex_ctrl_wb_sel~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_wb_sel~16 (
	.dataa(\ex_ctrl_wb_sel~15_combout ),
	.datab(\ex_ctrl_wb_sel~10_combout ),
	.datac(\ex_ctrl_wb_sel~12_combout ),
	.datad(\Equal50~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_wb_sel~16_combout ),
	.cout());
defparam \ex_ctrl_wb_sel~16 .lut_mask = 16'h2AEA;
defparam \ex_ctrl_wb_sel~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_wb_sel~17 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\ex_ctrl_wb_sel~16_combout ),
	.datad(\Equal5~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_wb_sel~17_combout ),
	.cout());
defparam \ex_ctrl_wb_sel~17 .lut_mask = 16'h0080;
defparam \ex_ctrl_wb_sel~17 .sum_lutc_input = "datac";

dffeas \ex_ctrl_wb_sel.00 (
	.clk(clk_clk),
	.d(\ex_ctrl_wb_sel~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_wb_sel.00~q ),
	.prn(vcc));
defparam \ex_ctrl_wb_sel.00 .is_wysiwyg = "true";
defparam \ex_ctrl_wb_sel.00 .power_up = "low";

cyclone10lp_lcell_comb \mem_ctrl_wb_sel~12 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_ctrl_wb_sel.00~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_ctrl_wb_sel~12_combout ),
	.cout());
defparam \mem_ctrl_wb_sel~12 .lut_mask = 16'h8888;
defparam \mem_ctrl_wb_sel~12 .sum_lutc_input = "datac";

dffeas \mem_ctrl_wb_sel.00 (
	.clk(clk_clk),
	.d(\mem_ctrl_wb_sel~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_ctrl_wb_sel.00~q ),
	.prn(vcc));
defparam \mem_ctrl_wb_sel.00 .is_wysiwyg = "true";
defparam \mem_ctrl_wb_sel.00 .power_up = "low";

cyclone10lp_lcell_comb \wb_ctrl_wb_sel~12 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_ctrl_wb_sel.00~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_ctrl_wb_sel~12_combout ),
	.cout());
defparam \wb_ctrl_wb_sel~12 .lut_mask = 16'h8888;
defparam \wb_ctrl_wb_sel~12 .sum_lutc_input = "datac";

dffeas \wb_ctrl_wb_sel.00 (
	.clk(clk_clk),
	.d(\wb_ctrl_wb_sel~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_ctrl_wb_sel.00~q ),
	.prn(vcc));
defparam \wb_ctrl_wb_sel.00 .is_wysiwyg = "true";
defparam \wb_ctrl_wb_sel.00 .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[23]~1 (
	.dataa(\wb_ctrl_wb_sel.10~q ),
	.datab(\wb_ctrl_wb_sel.00~q ),
	.datac(gnd),
	.datad(\wb_ctrl_wb_sel.11~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[23]~1_combout ),
	.cout());
defparam \_T_3543__T_3854_data[23]~1 .lut_mask = 16'hAAEE;
defparam \_T_3543__T_3854_data[23]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_alu_out~18 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~18_combout ),
	.cout());
defparam \wb_alu_out~18 .lut_mask = 16'h8888;
defparam \wb_alu_out~18 .sum_lutc_input = "datac";

dffeas \wb_alu_out[4] (
	.clk(clk_clk),
	.d(\wb_alu_out~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[4]~q ),
	.prn(vcc));
defparam \wb_alu_out[4] .is_wysiwyg = "true";
defparam \wb_alu_out[4] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[4]~39 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[4]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[4]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[4]~39_combout ),
	.cout());
defparam \_T_3543__T_3854_data[4]~39 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[4]~39 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~60 (
	.dataa(av_readdata_pre_28),
	.datab(av_readdata_pre_12),
	.datac(gnd),
	.datad(mem_alu_out_1),
	.cin(gnd),
	.combout(\wb_dmem_read_data~60_combout ),
	.cout());
defparam \wb_dmem_read_data~60 .lut_mask = 16'hAACC;
defparam \wb_dmem_read_data~60 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mask_type~4 (
	.dataa(\Equal15~1_combout ),
	.datab(\Equal8~1_combout ),
	.datac(\Equal17~0_combout ),
	.datad(\Equal18~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_mask_type~4_combout ),
	.cout());
defparam \ex_ctrl_mask_type~4 .lut_mask = 16'hEEEA;
defparam \ex_ctrl_mask_type~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mask_type~5 (
	.dataa(\ex_ctrl_mask_type~4_combout ),
	.datab(\Equal20~0_combout ),
	.datac(\ex_ctrl_mask_type~3_combout ),
	.datad(\Equal5~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_mask_type~5_combout ),
	.cout());
defparam \ex_ctrl_mask_type~5 .lut_mask = 16'hAAEA;
defparam \ex_ctrl_mask_type~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mask_type~6 (
	.dataa(\ex_ctrl_mem_wr~9_combout ),
	.datab(\id_pc[7]~31_combout ),
	.datac(\ex_ctrl_mask_type~5_combout ),
	.datad(\ex_ctrl_mem_wr~8_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_mask_type~6_combout ),
	.cout());
defparam \ex_ctrl_mask_type~6 .lut_mask = 16'hAABA;
defparam \ex_ctrl_mask_type~6 .sum_lutc_input = "datac";

dffeas \ex_ctrl_mask_type[0] (
	.clk(clk_clk),
	.d(\ex_ctrl_mask_type~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_mask_type[0]~q ),
	.prn(vcc));
defparam \ex_ctrl_mask_type[0] .is_wysiwyg = "true";
defparam \ex_ctrl_mask_type[0] .power_up = "low";

cyclone10lp_lcell_comb \mem_ctrl_mask_type~0 (
	.dataa(\ex_ctrl_mask_type[0]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_ctrl_mask_type~0_combout ),
	.cout());
defparam \mem_ctrl_mask_type~0 .lut_mask = 16'h8888;
defparam \mem_ctrl_mask_type~0 .sum_lutc_input = "datac";

dffeas \mem_ctrl_mask_type[0] (
	.clk(clk_clk),
	.d(\mem_ctrl_mask_type~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_ctrl_mask_type[0]~q ),
	.prn(vcc));
defparam \mem_ctrl_mask_type[0] .is_wysiwyg = "true";
defparam \mem_ctrl_mask_type[0] .power_up = "low";

cyclone10lp_lcell_comb \ex_ctrl_mask_type~8 (
	.dataa(\id_inst[12]~q ),
	.datab(\Equal18~1_combout ),
	.datac(\id_inst[4]~q ),
	.datad(\ex_ctrl_mask_type~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_mask_type~8_combout ),
	.cout());
defparam \ex_ctrl_mask_type~8 .lut_mask = 16'h08FF;
defparam \ex_ctrl_mask_type~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mask_type~9 (
	.dataa(\ex_ctrl_mask_type~8_combout ),
	.datab(\ex_ctrl_mask_type~3_combout ),
	.datac(\Equal5~1_combout ),
	.datad(\Equal20~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_mask_type~9_combout ),
	.cout());
defparam \ex_ctrl_mask_type~9 .lut_mask = 16'hAAAE;
defparam \ex_ctrl_mask_type~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mask_type~10 (
	.dataa(\ex_ctrl_mem_wr~9_combout ),
	.datab(\id_pc[7]~31_combout ),
	.datac(\ex_ctrl_mask_type~9_combout ),
	.datad(\ex_ctrl_mem_wr~8_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_mask_type~10_combout ),
	.cout());
defparam \ex_ctrl_mask_type~10 .lut_mask = 16'hAABA;
defparam \ex_ctrl_mask_type~10 .sum_lutc_input = "datac";

dffeas \ex_ctrl_mask_type[1] (
	.clk(clk_clk),
	.d(\ex_ctrl_mask_type~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_mask_type[1]~q ),
	.prn(vcc));
defparam \ex_ctrl_mask_type[1] .is_wysiwyg = "true";
defparam \ex_ctrl_mask_type[1] .power_up = "low";

cyclone10lp_lcell_comb \mem_ctrl_mask_type~2 (
	.dataa(\ex_ctrl_mask_type[1]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_ctrl_mask_type~2_combout ),
	.cout());
defparam \mem_ctrl_mask_type~2 .lut_mask = 16'h8888;
defparam \mem_ctrl_mask_type~2 .sum_lutc_input = "datac";

dffeas \mem_ctrl_mask_type[1] (
	.clk(clk_clk),
	.d(\mem_ctrl_mask_type~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_ctrl_mask_type[1]~q ),
	.prn(vcc));
defparam \mem_ctrl_mask_type[1] .is_wysiwyg = "true";
defparam \mem_ctrl_mask_type[1] .power_up = "low";

cyclone10lp_lcell_comb \wb_dmem_read_data[7]~17 (
	.dataa(mem_alu_out_1),
	.datab(\mem_ctrl_mask_type[0]~q ),
	.datac(\mem_ctrl_mask_type[1]~q ),
	.datad(mem_alu_out_0),
	.cin(gnd),
	.combout(\wb_dmem_read_data[7]~17_combout ),
	.cout());
defparam \wb_dmem_read_data[7]~17 .lut_mask = 16'h0028;
defparam \wb_dmem_read_data[7]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[4]~4 (
	.dataa(\wb_dmem_read_data~60_combout ),
	.datab(av_readdata_pre_20),
	.datac(gnd),
	.datad(\wb_dmem_read_data[7]~17_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data[4]~4_combout ),
	.cout());
defparam \wb_dmem_read_data[4]~4 .lut_mask = 16'hCCAA;
defparam \wb_dmem_read_data[4]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[7]~18 (
	.dataa(mem_alu_out_0),
	.datab(\mem_ctrl_mask_type[1]~q ),
	.datac(mem_ctrl_mem_wr01),
	.datad(\mem_ctrl_mask_type[0]~q ),
	.cin(gnd),
	.combout(\wb_dmem_read_data[7]~18_combout ),
	.cout());
defparam \wb_dmem_read_data[7]~18 .lut_mask = 16'h0080;
defparam \wb_dmem_read_data[7]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[7]~19 (
	.dataa(\wb_dmem_read_data[7]~18_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\wb_dmem_read_data[7]~19_combout ),
	.cout());
defparam \wb_dmem_read_data[7]~19 .lut_mask = 16'hAAFF;
defparam \wb_dmem_read_data[7]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[7]~20 (
	.dataa(\mem_ctrl_mask_type[0]~q ),
	.datab(\mem_ctrl_mask_type[1]~q ),
	.datac(mem_alu_out_0),
	.datad(mem_alu_out_1),
	.cin(gnd),
	.combout(\wb_dmem_read_data[7]~20_combout ),
	.cout());
defparam \wb_dmem_read_data[7]~20 .lut_mask = 16'h999F;
defparam \wb_dmem_read_data[7]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[7]~21 (
	.dataa(\wb_dmem_read_data[7]~20_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_ctrl_mem_wr01),
	.cin(gnd),
	.combout(\wb_dmem_read_data[7]~21_combout ),
	.cout());
defparam \wb_dmem_read_data[7]~21 .lut_mask = 16'hAAFF;
defparam \wb_dmem_read_data[7]~21 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[4] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data[4]~4_combout ),
	.asdata(av_readdata_pre_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\wb_dmem_read_data[7]~19_combout ),
	.sload(\wb_dmem_read_data[7]~21_combout ),
	.ena(vcc),
	.q(\wb_dmem_read_data[4]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[4] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[4] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[4]~40 (
	.dataa(\wb_csr_data[4]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[4]~39_combout ),
	.datad(\wb_dmem_read_data[4]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[4]~40_combout ),
	.cout());
defparam \_T_3543__T_3854_data[4]~40 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[4]~40 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a28 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[4]~40_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a28_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_a_first_bit_number = 28;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_b_first_bit_number = 28;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a28 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~20 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a28~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~20_combout ),
	.cout());
defparam \ex_rs_1~20 .lut_mask = 16'h8888;
defparam \ex_rs_1~20 .sum_lutc_input = "datac";

dffeas \ex_rs_1[4] (
	.clk(clk_clk),
	.d(\ex_rs_1~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[4]~q ),
	.prn(vcc));
defparam \ex_rs_1[4] .is_wysiwyg = "true";
defparam \ex_rs_1[4] .power_up = "low";

cyclone10lp_lcell_comb \wb_ctrl_csr_cmd~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\mem_ctrl_csr_cmd.000~q ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\wb_ctrl_csr_cmd~14_combout ),
	.cout());
defparam \wb_ctrl_csr_cmd~14 .lut_mask = 16'hF000;
defparam \wb_ctrl_csr_cmd~14 .sum_lutc_input = "datac";

dffeas \wb_ctrl_csr_cmd.000 (
	.clk(clk_clk),
	.d(\wb_ctrl_csr_cmd~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_ctrl_csr_cmd.000~q ),
	.prn(vcc));
defparam \wb_ctrl_csr_cmd.000 .is_wysiwyg = "true";
defparam \wb_ctrl_csr_cmd.000 .power_up = "low";

cyclone10lp_lcell_comb \Equal53~1 (
	.dataa(\Equal53~0_combout ),
	.datab(\Equal18~0_combout ),
	.datac(gnd),
	.datad(\id_inst[14]~q ),
	.cin(gnd),
	.combout(\Equal53~1_combout ),
	.cout());
defparam \Equal53~1 .lut_mask = 16'h0088;
defparam \Equal53~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb _T_3091(
	.dataa(\Equal8~1_combout ),
	.datab(\_T_3083~0_combout ),
	.datac(\Equal53~1_combout ),
	.datad(\_T_3091~0_combout ),
	.cin(gnd),
	.combout(\_T_3091~combout ),
	.cout());
defparam _T_3091.lut_mask = 16'h80FF;
defparam _T_3091.sum_lutc_input = "datac";

cyclone10lp_lcell_comb _GEN_15(
	.dataa(\_T_1778~combout ),
	.datab(\_GEN_15~2_combout ),
	.datac(\_T_3091~combout ),
	.datad(\Equal5~1_combout ),
	.cin(gnd),
	.combout(\_GEN_15~combout ),
	.cout());
defparam _GEN_15.lut_mask = 16'h0080;
defparam _GEN_15.sum_lutc_input = "datac";

dffeas ex_ctrl_mem_en(
	.clk(clk_clk),
	.d(\_GEN_15~combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_mem_en~q ),
	.prn(vcc));
defparam ex_ctrl_mem_en.is_wysiwyg = "true";
defparam ex_ctrl_mem_en.power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[2]~8 (
	.dataa(\ex_ctrl_rf_wen~q ),
	.datab(\wb_ctrl_csr_cmd.000~q ),
	.datac(\wb_ctrl_rf_wen~q ),
	.datad(\ex_ctrl_mem_en~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[2]~8_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[2]~8 .lut_mask = 16'h8ACF;
defparam \ex_reg_rs1_bypass[2]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal64~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\ex_csr_addr[4]~q ),
	.datad(\wb_reg_waddr[4]~q ),
	.cin(gnd),
	.combout(\Equal64~0_combout ),
	.cout());
defparam \Equal64~0 .lut_mask = 16'h0FF0;
defparam \Equal64~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3689~0 (
	.dataa(\ex_csr_addr[0]~q ),
	.datab(\ex_csr_addr[1]~q ),
	.datac(\wb_reg_waddr[1]~q ),
	.datad(\wb_reg_waddr[0]~q ),
	.cin(gnd),
	.combout(\_T_3689~0_combout ),
	.cout());
defparam \_T_3689~0 .lut_mask = 16'h8241;
defparam \_T_3689~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3689~1 (
	.dataa(\ex_csr_addr[2]~q ),
	.datab(\wb_reg_waddr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\_T_3689~1_combout ),
	.cout());
defparam \_T_3689~1 .lut_mask = 16'h9999;
defparam \_T_3689~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3689~2 (
	.dataa(\ex_csr_addr[3]~q ),
	.datab(\wb_reg_waddr[3]~q ),
	.datac(\_T_3689~0_combout ),
	.datad(\_T_3689~1_combout ),
	.cin(gnd),
	.combout(\_T_3689~2_combout ),
	.cout());
defparam \_T_3689~2 .lut_mask = 16'h9000;
defparam \_T_3689~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[7]~4 (
	.dataa(\Equal62~1_combout ),
	.datab(\ex_reg_rs1_bypass[2]~8_combout ),
	.datac(\Equal64~0_combout ),
	.datad(\_T_3689~2_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[7]~4_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[7]~4 .lut_mask = 16'hFEFF;
defparam \ex_reg_rs2_bypass[7]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb _GEN_39(
	.dataa(\ex_ctrl_mem_en~q ),
	.datab(\inst_kill~0_combout ),
	.datac(\csr|io_expt~0_combout ),
	.datad(\csr|isEcall~0_combout ),
	.cin(gnd),
	.combout(\_GEN_39~combout ),
	.cout());
defparam _GEN_39.lut_mask = 16'h0080;
defparam _GEN_39.sum_lutc_input = "datac";

dffeas mem_ctrl_mem_en(
	.clk(clk_clk),
	.d(\_GEN_39~combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_ctrl_mem_en~q ),
	.prn(vcc));
defparam mem_ctrl_mem_en.is_wysiwyg = "true";
defparam mem_ctrl_mem_en.power_up = "low";

cyclone10lp_lcell_comb \wb_ctrl_mem_en~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_ctrl_mem_en~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_ctrl_mem_en~0_combout ),
	.cout());
defparam \wb_ctrl_mem_en~0 .lut_mask = 16'h8888;
defparam \wb_ctrl_mem_en~0 .sum_lutc_input = "datac";

dffeas wb_ctrl_mem_en(
	.clk(clk_clk),
	.d(\wb_ctrl_mem_en~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_ctrl_mem_en~q ),
	.prn(vcc));
defparam wb_ctrl_mem_en.is_wysiwyg = "true";
defparam wb_ctrl_mem_en.power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[2]~6 (
	.dataa(\ex_ctrl_rf_wen~q ),
	.datab(\wb_ctrl_mem_en~q ),
	.datac(\wb_ctrl_csr_cmd.000~q ),
	.datad(\ex_ctrl_mem_en~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[2]~6_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[2]~6 .lut_mask = 16'hACFC;
defparam \ex_reg_rs1_bypass[2]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[2]~12 (
	.dataa(\wb_ctrl_rf_wen~q ),
	.datab(\ex_reg_rs1_bypass[2]~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[2]~12_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[2]~12 .lut_mask = 16'h8888;
defparam \ex_reg_rs1_bypass[2]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[7]~5 (
	.dataa(\_T_3689~2_combout ),
	.datab(\ex_reg_rs1_bypass[2]~12_combout ),
	.datac(\Equal62~1_combout ),
	.datad(\Equal64~0_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[7]~5_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[7]~5 .lut_mask = 16'h0008;
defparam \ex_reg_rs2_bypass[7]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[4]~75 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_4),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[4]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[4]~75_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[4]~75 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[4]~75 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[4]~76 (
	.dataa(\ex_rs_1[4]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[4]~75_combout ),
	.datad(\wb_csr_data[4]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[4]~76_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[4]~76 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[4]~76 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[4]~60 (
	.dataa(\mem_alu_out[4]~q ),
	.datab(\_T_3686~0_combout ),
	.datac(\ex_reg_rs2_bypass[4]~76_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\alu_io_op2[4]~60_combout ),
	.cout());
defparam \alu_io_op2[4]~60 .lut_mask = 16'hB8B8;
defparam \alu_io_op2[4]~60 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[4]~61 (
	.dataa(\ex_ctrl_alu_op2.10~q ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[4]~q ),
	.datad(\alu_io_op2[4]~60_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[4]~61_combout ),
	.cout());
defparam \alu_io_op2[4]~61 .lut_mask = 16'hA280;
defparam \alu_io_op2[4]~61 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[4]~62 (
	.dataa(\csr_io_alu_op2[1]~0_combout ),
	.datab(\alu_io_op2[4]~61_combout ),
	.datac(\io_sw_r_ex_imm[4]~4_combout ),
	.datad(\ex_ctrl_alu_op2.10~q ),
	.cin(gnd),
	.combout(\alu_io_op2[4]~62_combout ),
	.cout());
defparam \alu_io_op2[4]~62 .lut_mask = 16'h88A8;
defparam \alu_io_op2[4]~62 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~16 (
	.dataa(\Equal5~1_combout ),
	.datab(\ex_ctrl_csr_cmd~12_combout ),
	.datac(gnd),
	.datad(\ex_csr_cmd~4_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~16_combout ),
	.cout());
defparam \ex_ctrl_alu_func~16 .lut_mask = 16'hAAEE;
defparam \ex_ctrl_alu_func~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal35~0 (
	.dataa(\id_inst[13]~q ),
	.datab(\Equal32~0_combout ),
	.datac(gnd),
	.datad(\id_inst[30]~q ),
	.cin(gnd),
	.combout(\Equal35~0_combout ),
	.cout());
defparam \Equal35~0 .lut_mask = 16'h0088;
defparam \Equal35~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal36~0 (
	.dataa(\id_inst[12]~q ),
	.datab(\Equal35~0_combout ),
	.datac(gnd),
	.datad(\id_inst[14]~q ),
	.cin(gnd),
	.combout(\Equal36~0_combout ),
	.cout());
defparam \Equal36~0 .lut_mask = 16'h0088;
defparam \Equal36~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~17 (
	.dataa(\Equal36~0_combout ),
	.datab(\Equal37~0_combout ),
	.datac(\ex_ctrl_imm_type~13_combout ),
	.datad(\Equal34~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~17_combout ),
	.cout());
defparam \ex_ctrl_alu_func~17 .lut_mask = 16'h00BA;
defparam \ex_ctrl_alu_func~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~18 (
	.dataa(\Equal31~1_combout ),
	.datab(\Equal33~0_combout ),
	.datac(\ex_ctrl_alu_func~17_combout ),
	.datad(\Equal32~2_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~18_combout ),
	.cout());
defparam \ex_ctrl_alu_func~18 .lut_mask = 16'hAAFE;
defparam \ex_ctrl_alu_func~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~19 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\Equal28~1_combout ),
	.datad(\Equal27~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~19_combout ),
	.cout());
defparam \ex_ctrl_alu_func~19 .lut_mask = 16'h000F;
defparam \ex_ctrl_alu_func~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~20 (
	.dataa(\ex_ctrl_alu_func~5_combout ),
	.datab(\ex_ctrl_alu_func~18_combout ),
	.datac(\ex_ctrl_alu_func~19_combout ),
	.datad(\Equal26~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~20_combout ),
	.cout());
defparam \ex_ctrl_alu_func~20 .lut_mask = 16'h0080;
defparam \ex_ctrl_alu_func~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~21 (
	.dataa(\ex_ctrl_alu_func~9_combout ),
	.datab(\ex_ctrl_alu_func~20_combout ),
	.datac(\ex_ctrl_alu_func~6_combout ),
	.datad(\Equal11~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~21_combout ),
	.cout());
defparam \ex_ctrl_alu_func~21 .lut_mask = 16'hFF8A;
defparam \ex_ctrl_alu_func~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~22 (
	.dataa(\ex_ctrl_alu_func~4_combout ),
	.datab(\ex_ctrl_alu_op1~2_combout ),
	.datac(\Equal8~2_combout ),
	.datad(\ex_ctrl_csr_cmd~12_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~22_combout ),
	.cout());
defparam \ex_ctrl_alu_func~22 .lut_mask = 16'h0002;
defparam \ex_ctrl_alu_func~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~23 (
	.dataa(\id_pc[7]~31_combout ),
	.datab(\ex_ctrl_alu_func~16_combout ),
	.datac(\ex_ctrl_alu_func~21_combout ),
	.datad(\ex_ctrl_alu_func~22_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~23_combout ),
	.cout());
defparam \ex_ctrl_alu_func~23 .lut_mask = 16'h5444;
defparam \ex_ctrl_alu_func~23 .sum_lutc_input = "datac";

dffeas \ex_ctrl_alu_func[3] (
	.clk(clk_clk),
	.d(\ex_ctrl_alu_func~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_alu_func[3]~q ),
	.prn(vcc));
defparam \ex_ctrl_alu_func[3] .is_wysiwyg = "true";
defparam \ex_ctrl_alu_func[3] .power_up = "low";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~24 (
	.dataa(\ex_ctrl_alu_op1~2_combout ),
	.datab(\ex_ctrl_mask_type~0_combout ),
	.datac(gnd),
	.datad(\Equal8~2_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~24_combout ),
	.cout());
defparam \ex_ctrl_alu_func~24 .lut_mask = 16'h0044;
defparam \ex_ctrl_alu_func~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~25 (
	.dataa(\Equal31~1_combout ),
	.datab(\id_inst[13]~q ),
	.datac(\Equal37~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~25_combout ),
	.cout());
defparam \ex_ctrl_alu_func~25 .lut_mask = 16'hEAEA;
defparam \ex_ctrl_alu_func~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~26 (
	.dataa(\ex_ctrl_alu_func~5_combout ),
	.datab(\Equal36~0_combout ),
	.datac(\ex_ctrl_alu_func~25_combout ),
	.datad(\ex_ctrl_alu_func~8_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~26_combout ),
	.cout());
defparam \ex_ctrl_alu_func~26 .lut_mask = 16'hA8AA;
defparam \ex_ctrl_alu_func~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~27 (
	.dataa(\Equal28~1_combout ),
	.datab(\Equal27~0_combout ),
	.datac(\ex_ctrl_alu_func~26_combout ),
	.datad(\Equal26~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~27_combout ),
	.cout());
defparam \ex_ctrl_alu_func~27 .lut_mask = 16'h00FE;
defparam \ex_ctrl_alu_func~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~35 (
	.dataa(\Equal17~0_combout ),
	.datab(\id_inst[4]~q ),
	.datac(\ex_ctrl_alu_func~27_combout ),
	.datad(\id_inst[12]~q ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~35_combout ),
	.cout());
defparam \ex_ctrl_alu_func~35 .lut_mask = 16'hF870;
defparam \ex_ctrl_alu_func~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~36 (
	.dataa(\ex_ctrl_alu_func~9_combout ),
	.datab(\ex_ctrl_alu_func~35_combout ),
	.datac(\Equal11~0_combout ),
	.datad(\id_inst[13]~q ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~36_combout ),
	.cout());
defparam \ex_ctrl_alu_func~36 .lut_mask = 16'hF808;
defparam \ex_ctrl_alu_func~36 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~28 (
	.dataa(\ex_ctrl_alu_func~24_combout ),
	.datab(\ex_ctrl_alu_func~36_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_func~4_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~28_combout ),
	.cout());
defparam \ex_ctrl_alu_func~28 .lut_mask = 16'h88AA;
defparam \ex_ctrl_alu_func~28 .sum_lutc_input = "datac";

dffeas \ex_ctrl_alu_func[1] (
	.clk(clk_clk),
	.d(\ex_ctrl_alu_func~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_alu_func[1]~q ),
	.prn(vcc));
defparam \ex_ctrl_alu_func[1] .is_wysiwyg = "true";
defparam \ex_ctrl_alu_func[1] .power_up = "low";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~29 (
	.dataa(\id_inst[14]~q ),
	.datab(\Equal29~1_combout ),
	.datac(\Equal31~1_combout ),
	.datad(\ex_csr_cmd~10_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~29_combout ),
	.cout());
defparam \ex_ctrl_alu_func~29 .lut_mask = 16'h888F;
defparam \ex_ctrl_alu_func~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~30 (
	.dataa(\ex_ctrl_alu_func~29_combout ),
	.datab(\id_inst[14]~q ),
	.datac(\id_inst[25]~q ),
	.datad(\Equal29~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~30_combout ),
	.cout());
defparam \ex_ctrl_alu_func~30 .lut_mask = 16'hA8AA;
defparam \ex_ctrl_alu_func~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~31 (
	.dataa(\ex_ctrl_alu_func~9_combout ),
	.datab(\ex_ctrl_alu_func~30_combout ),
	.datac(\ex_ctrl_alu_func~7_combout ),
	.datad(\Equal11~0_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~31_combout ),
	.cout());
defparam \ex_ctrl_alu_func~31 .lut_mask = 16'hFF8A;
defparam \ex_ctrl_alu_func~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_func~32 (
	.dataa(\ex_ctrl_alu_func~4_combout ),
	.datab(\ex_ctrl_alu_func~24_combout ),
	.datac(\ex_ctrl_alu_func~31_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_ctrl_alu_func~32_combout ),
	.cout());
defparam \ex_ctrl_alu_func~32 .lut_mask = 16'h8080;
defparam \ex_ctrl_alu_func~32 .sum_lutc_input = "datac";

dffeas \ex_ctrl_alu_func[2] (
	.clk(clk_clk),
	.d(\ex_ctrl_alu_func~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_alu_func[2]~q ),
	.prn(vcc));
defparam \ex_ctrl_alu_func[2] .is_wysiwyg = "true";
defparam \ex_ctrl_alu_func[2] .power_up = "low";

cyclone10lp_lcell_comb \mem_alu_out[26]~0 (
	.dataa(\ex_ctrl_alu_func[0]~q ),
	.datab(\ex_ctrl_alu_func[3]~q ),
	.datac(\ex_ctrl_alu_func[1]~q ),
	.datad(\ex_ctrl_alu_func[2]~q ),
	.cin(gnd),
	.combout(\mem_alu_out[26]~0_combout ),
	.cout());
defparam \mem_alu_out[26]~0 .lut_mask = 16'h8AF8;
defparam \mem_alu_out[26]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_alu_op1~6 (
	.dataa(\ex_ctrl_alu_func~4_combout ),
	.datab(\Equal11~0_combout ),
	.datac(\ex_ctrl_imm_type~12_combout ),
	.datad(\ex_ctrl_alu_op1~5_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_alu_op1~6_combout ),
	.cout());
defparam \ex_ctrl_alu_op1~6 .lut_mask = 16'hDFFF;
defparam \ex_ctrl_alu_op1~6 .sum_lutc_input = "datac";

dffeas \ex_ctrl_alu_op1[0] (
	.clk(clk_clk),
	.d(\ex_ctrl_alu_op1~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!altera_reset_synchronizer_int_chain_out),
	.ena(vcc),
	.q(\ex_ctrl_alu_op1[0]~q ),
	.prn(vcc));
defparam \ex_ctrl_alu_op1[0] .is_wysiwyg = "true";
defparam \ex_ctrl_alu_op1[0] .power_up = "low";

dffeas \ex_ctrl_alu_op1[1] (
	.clk(clk_clk),
	.d(\ex_ctrl_alu_op1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\id_pc[7]~31_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_alu_op1[1]~q ),
	.prn(vcc));
defparam \ex_ctrl_alu_op1[1] .is_wysiwyg = "true";
defparam \ex_ctrl_alu_op1[1] .power_up = "low";

cyclone10lp_lcell_comb \Equal59~0 (
	.dataa(\ex_inst[15]~q ),
	.datab(\ex_inst[16]~q ),
	.datac(\ex_inst[17]~q ),
	.datad(\ex_inst[18]~q ),
	.cin(gnd),
	.combout(\Equal59~0_combout ),
	.cout());
defparam \Equal59~0 .lut_mask = 16'h0001;
defparam \Equal59~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal59~1 (
	.dataa(\Equal59~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ex_inst[19]~q ),
	.cin(gnd),
	.combout(\Equal59~1_combout ),
	.cout());
defparam \Equal59~1 .lut_mask = 16'h00AA;
defparam \Equal59~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal60~2 (
	.dataa(\mem_reg_waddr[0]~q ),
	.datab(\mem_reg_waddr[1]~q ),
	.datac(\ex_inst[16]~q ),
	.datad(\ex_inst[15]~q ),
	.cin(gnd),
	.combout(\Equal60~2_combout ),
	.cout());
defparam \Equal60~2 .lut_mask = 16'h8241;
defparam \Equal60~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal60~3 (
	.dataa(\mem_reg_waddr[2]~q ),
	.datab(\mem_reg_waddr[3]~q ),
	.datac(\ex_inst[18]~q ),
	.datad(\ex_inst[17]~q ),
	.cin(gnd),
	.combout(\Equal60~3_combout ),
	.cout());
defparam \Equal60~3 .lut_mask = 16'h8241;
defparam \Equal60~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal60~5 (
	.dataa(\mem_reg_waddr[4]~q ),
	.datab(\ex_inst[19]~q ),
	.datac(\Equal60~2_combout ),
	.datad(\Equal60~3_combout ),
	.cin(gnd),
	.combout(\Equal60~5_combout ),
	.cout());
defparam \Equal60~5 .lut_mask = 16'h9000;
defparam \Equal60~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal60~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\mem_reg_waddr[4]~q ),
	.datad(\ex_inst[19]~q ),
	.cin(gnd),
	.combout(\Equal60~4_combout ),
	.cout());
defparam \Equal60~4 .lut_mask = 16'h0FF0;
defparam \Equal60~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_in[0]~0 (
	.dataa(\mem_ctrl_csr_cmd.000~q ),
	.datab(\Equal60~2_combout ),
	.datac(\Equal60~3_combout ),
	.datad(\Equal60~4_combout ),
	.cin(gnd),
	.combout(\csr_io_in[0]~0_combout ),
	.cout());
defparam \csr_io_in[0]~0 .lut_mask = 16'h0080;
defparam \csr_io_in[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[0]~4 (
	.dataa(\Equal59~1_combout ),
	.datab(\mem_ctrl_rf_wen~q ),
	.datac(\Equal60~5_combout ),
	.datad(\csr_io_in[0]~0_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[0]~4_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[0]~4 .lut_mask = 16'hAABF;
defparam \ex_reg_rs1_bypass[0]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[0]~20 (
	.dataa(\mem_ctrl_rf_wen~q ),
	.datab(\Equal60~5_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\Equal59~1_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[0]~20_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[0]~20 .lut_mask = 16'h0008;
defparam \ex_reg_rs1_bypass[0]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3634~2 (
	.dataa(\Equal59~0_combout ),
	.datab(\ex_inst[19]~q ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\_T_3634~2_combout ),
	.cout());
defparam \_T_3634~2 .lut_mask = 16'hD0D0;
defparam \_T_3634~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[4]~82 (
	.dataa(\ex_reg_rs1_bypass[0]~20_combout ),
	.datab(\mem_alu_out[4]~q ),
	.datac(\_T_3634~2_combout ),
	.datad(\mem_csr_data[4]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[4]~82_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[4]~82 .lut_mask = 16'hF888;
defparam \ex_reg_rs1_bypass[4]~82 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a28 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[4]~40_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a28_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_a_first_bit_number = 28;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_b_first_bit_number = 28;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a28 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~20 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a28~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~20_combout ),
	.cout());
defparam \ex_rs_0~20 .lut_mask = 16'h0080;
defparam \ex_rs_0~20 .sum_lutc_input = "datac";

dffeas \ex_rs_0[4] (
	.clk(clk_clk),
	.d(\ex_rs_0~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[4]~q ),
	.prn(vcc));
defparam \ex_rs_0[4] .is_wysiwyg = "true";
defparam \ex_rs_0[4] .power_up = "low";

cyclone10lp_lcell_comb \Equal61~0 (
	.dataa(\wb_reg_waddr[0]~q ),
	.datab(\wb_reg_waddr[1]~q ),
	.datac(\ex_inst[16]~q ),
	.datad(\ex_inst[15]~q ),
	.cin(gnd),
	.combout(\Equal61~0_combout ),
	.cout());
defparam \Equal61~0 .lut_mask = 16'h8241;
defparam \Equal61~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal61~1 (
	.dataa(\wb_reg_waddr[2]~q ),
	.datab(\wb_reg_waddr[3]~q ),
	.datac(\ex_inst[18]~q ),
	.datad(\ex_inst[17]~q ),
	.cin(gnd),
	.combout(\Equal61~1_combout ),
	.cout());
defparam \Equal61~1 .lut_mask = 16'h8241;
defparam \Equal61~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal61~2 (
	.dataa(\Equal61~0_combout ),
	.datab(\Equal61~1_combout ),
	.datac(\wb_reg_waddr[4]~q ),
	.datad(\ex_inst[19]~q ),
	.cin(gnd),
	.combout(\Equal61~2_combout ),
	.cout());
defparam \Equal61~2 .lut_mask = 16'h8008;
defparam \Equal61~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[2]~138 (
	.dataa(\Equal59~0_combout ),
	.datab(\ex_inst[19]~q ),
	.datac(\ex_reg_rs1_bypass[2]~8_combout ),
	.datad(\Equal61~2_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[2]~138_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[2]~138 .lut_mask = 16'hF2FF;
defparam \ex_reg_rs1_bypass[2]~138 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[2]~7 (
	.dataa(\wb_ctrl_rf_wen~q ),
	.datab(\ex_reg_rs1_bypass[2]~6_combout ),
	.datac(\Equal61~2_combout ),
	.datad(\Equal59~1_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[2]~7_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[2]~7 .lut_mask = 16'h0080;
defparam \ex_reg_rs1_bypass[2]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[4]~83 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(av_readdata_pre_4),
	.datac(\wb_alu_out[4]~q ),
	.datad(\ex_reg_rs1_bypass[2]~138_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[4]~83_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[4]~83 .lut_mask = 16'hAAD8;
defparam \ex_reg_rs1_bypass[4]~83 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[4]~84 (
	.dataa(\ex_rs_0[4]~q ),
	.datab(\wb_csr_data[4]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\ex_reg_rs1_bypass[4]~83_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[4]~84_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[4]~84 .lut_mask = 16'hCFA0;
defparam \ex_reg_rs1_bypass[4]~84 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[4]~85 (
	.dataa(\ex_reg_rs1_bypass[0]~4_combout ),
	.datab(\ex_reg_rs1_bypass[4]~82_combout ),
	.datac(\ex_reg_rs1_bypass[4]~84_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[4]~85_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[4]~85 .lut_mask = 16'hECEC;
defparam \ex_reg_rs1_bypass[4]~85 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[4]~106 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[4]~q ),
	.datad(\ex_reg_rs1_bypass[4]~85_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[4]~106_combout ),
	.cout());
defparam \alu_io_op1[4]~106 .lut_mask = 16'h6240;
defparam \alu_io_op1[4]~106 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out[26]~1 (
	.dataa(\ex_ctrl_alu_func[3]~q ),
	.datab(\ex_ctrl_alu_func[1]~q ),
	.datac(\ex_ctrl_alu_func[2]~q ),
	.datad(\ex_ctrl_alu_func[0]~q ),
	.cin(gnd),
	.combout(\mem_alu_out[26]~1_combout ),
	.cout());
defparam \mem_alu_out[26]~1 .lut_mask = 16'h18AA;
defparam \mem_alu_out[26]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out[26]~2 (
	.dataa(\ex_ctrl_alu_func[2]~q ),
	.datab(\ex_ctrl_alu_func[0]~q ),
	.datac(gnd),
	.datad(\ex_ctrl_alu_func[1]~q ),
	.cin(gnd),
	.combout(\mem_alu_out[26]~2_combout ),
	.cout());
defparam \mem_alu_out[26]~2 .lut_mask = 16'h88AA;
defparam \mem_alu_out[26]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~143 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\alu_io_op2[4]~62_combout ),
	.datad(\alu_io_op1[4]~106_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~143_combout ),
	.cout());
defparam \mem_alu_out~143 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~143 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~144 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~143_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~251_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~144_combout ),
	.cout());
defparam \mem_alu_out~144 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~144 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~85 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[4]~106_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~144_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~85_combout ),
	.cout());
defparam \mem_alu_out~85 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~85 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~86 (
	.dataa(\alu_io_op2[4]~62_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~85_combout ),
	.datad(\alu|ShiftRight0~228_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~86_combout ),
	.cout());
defparam \mem_alu_out~86 .lut_mask = 16'hF838;
defparam \mem_alu_out~86 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out[26]~5 (
	.dataa(\ex_ctrl_alu_func[0]~q ),
	.datab(\ex_ctrl_alu_func[2]~q ),
	.datac(\ex_ctrl_alu_func[3]~q ),
	.datad(\ex_ctrl_alu_func[1]~q ),
	.cin(gnd),
	.combout(\mem_alu_out[26]~5_combout ),
	.cout());
defparam \mem_alu_out[26]~5 .lut_mask = 16'hEFFE;
defparam \mem_alu_out[26]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out[26]~6 (
	.dataa(\ex_ctrl_alu_func[3]~q ),
	.datab(\ex_ctrl_alu_func[2]~q ),
	.datac(\ex_ctrl_alu_func[0]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_alu_out[26]~6_combout ),
	.cout());
defparam \mem_alu_out[26]~6 .lut_mask = 16'h08FF;
defparam \mem_alu_out[26]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~87 (
	.dataa(\mem_alu_out~86_combout ),
	.datab(\alu|_T_3[4]~8_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~87_combout ),
	.cout());
defparam \mem_alu_out~87 .lut_mask = 16'h00AC;
defparam \mem_alu_out~87 .sum_lutc_input = "datac";

dffeas \mem_alu_out[4] (
	.clk(clk_clk),
	.d(\mem_alu_out~87_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[4]~q ),
	.prn(vcc));
defparam \mem_alu_out[4] .is_wysiwyg = "true";
defparam \mem_alu_out[4] .power_up = "low";

cyclone10lp_lcell_comb \pc_cntr~16 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(\mem_alu_out[4]~q ),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[4]~4_combout ),
	.cin(gnd),
	.combout(\pc_cntr~16_combout ),
	.cout());
defparam \pc_cntr~16 .lut_mask = 16'hDAD0;
defparam \pc_cntr~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~17 (
	.dataa(\_T_3862[4]~8_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~16_combout ),
	.datad(\csr|mepc[4]~q ),
	.cin(gnd),
	.combout(\pc_cntr~17_combout ),
	.cout());
defparam \pc_cntr~17 .lut_mask = 16'hF2C2;
defparam \pc_cntr~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~18 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~17_combout ),
	.datac(\csr|mtvec[4]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~18_combout ),
	.cout());
defparam \pc_cntr~18 .lut_mask = 16'h88A0;
defparam \pc_cntr~18 .sum_lutc_input = "datac";

dffeas \pc_cntr[4] (
	.clk(clk_clk),
	.d(\pc_cntr~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[4]~q ),
	.prn(vcc));
defparam \pc_cntr[4] .is_wysiwyg = "true";
defparam \pc_cntr[4] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~3 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~3_combout ),
	.cout());
defparam \id_pc~3 .lut_mask = 16'h8080;
defparam \id_pc~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~1 (
	.dataa(id_pc_5),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~1_combout ),
	.cout());
defparam \ex_pc~1 .lut_mask = 16'h8080;
defparam \ex_pc~1 .sum_lutc_input = "datac";

dffeas \ex_pc[5] (
	.clk(clk_clk),
	.d(\ex_pc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[5]~q ),
	.prn(vcc));
defparam \ex_pc[5] .is_wysiwyg = "true";
defparam \ex_pc[5] .power_up = "low";

cyclone10lp_lcell_comb \mem_csr_data~28 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[5]~166_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~28_combout ),
	.cout());
defparam \mem_csr_data~28 .lut_mask = 16'h8888;
defparam \mem_csr_data~28 .sum_lutc_input = "datac";

dffeas \mem_csr_data[5] (
	.clk(clk_clk),
	.d(\mem_csr_data~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[5]~q ),
	.prn(vcc));
defparam \mem_csr_data[5] .is_wysiwyg = "true";
defparam \mem_csr_data[5] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[5]~90 (
	.dataa(\ex_reg_rs1_bypass[0]~20_combout ),
	.datab(\mem_alu_out[5]~q ),
	.datac(\_T_3634~2_combout ),
	.datad(\mem_csr_data[5]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[5]~90_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[5]~90 .lut_mask = 16'hF888;
defparam \ex_reg_rs1_bypass[5]~90 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_csr_data~21 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~21_combout ),
	.cout());
defparam \wb_csr_data~21 .lut_mask = 16'h8888;
defparam \wb_csr_data~21 .sum_lutc_input = "datac";

dffeas \wb_csr_data[5] (
	.clk(clk_clk),
	.d(\wb_csr_data~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[5]~q ),
	.prn(vcc));
defparam \wb_csr_data[5] .is_wysiwyg = "true";
defparam \wb_csr_data[5] .power_up = "low";

cyclone10lp_lcell_comb \npc[5]~6 (
	.dataa(\pc_cntr[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[4]~5 ),
	.combout(\npc[5]~6_combout ),
	.cout(\npc[5]~7 ));
defparam \npc[5]~6 .lut_mask = 16'h5A5F;
defparam \npc[5]~6 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~21 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[5]~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~21_combout ),
	.cout());
defparam \id_npc~21 .lut_mask = 16'h8080;
defparam \id_npc~21 .sum_lutc_input = "datac";

dffeas \id_npc[5] (
	.clk(clk_clk),
	.d(\id_npc~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[5]~q ),
	.prn(vcc));
defparam \id_npc[5] .is_wysiwyg = "true";
defparam \id_npc[5] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~21 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~21_combout ),
	.cout());
defparam \ex_npc~21 .lut_mask = 16'h8080;
defparam \ex_npc~21 .sum_lutc_input = "datac";

dffeas \ex_npc[5] (
	.clk(clk_clk),
	.d(\ex_npc~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[5]~q ),
	.prn(vcc));
defparam \ex_npc[5] .is_wysiwyg = "true";
defparam \ex_npc[5] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~19 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~19_combout ),
	.cout());
defparam \mem_npc~19 .lut_mask = 16'h8888;
defparam \mem_npc~19 .sum_lutc_input = "datac";

dffeas \mem_npc[5] (
	.clk(clk_clk),
	.d(\mem_npc~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[5]~q ),
	.prn(vcc));
defparam \mem_npc[5] .is_wysiwyg = "true";
defparam \mem_npc[5] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~19 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~19_combout ),
	.cout());
defparam \wb_npc~19 .lut_mask = 16'h8888;
defparam \wb_npc~19 .sum_lutc_input = "datac";

dffeas \wb_npc[5] (
	.clk(clk_clk),
	.d(\wb_npc~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[5]~q ),
	.prn(vcc));
defparam \wb_npc[5] .is_wysiwyg = "true";
defparam \wb_npc[5] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~21 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~21_combout ),
	.cout());
defparam \wb_alu_out~21 .lut_mask = 16'h8888;
defparam \wb_alu_out~21 .sum_lutc_input = "datac";

dffeas \wb_alu_out[5] (
	.clk(clk_clk),
	.d(\wb_alu_out~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[5]~q ),
	.prn(vcc));
defparam \wb_alu_out[5] .is_wysiwyg = "true";
defparam \wb_alu_out[5] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[5]~45 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[5]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[5]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[5]~45_combout ),
	.cout());
defparam \_T_3543__T_3854_data[5]~45 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[5]~45 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~64 (
	.dataa(av_readdata_pre_29),
	.datab(av_readdata_pre_13),
	.datac(gnd),
	.datad(mem_alu_out_1),
	.cin(gnd),
	.combout(\wb_dmem_read_data~64_combout ),
	.cout());
defparam \wb_dmem_read_data~64 .lut_mask = 16'hAACC;
defparam \wb_dmem_read_data~64 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[5]~3 (
	.dataa(\wb_dmem_read_data~64_combout ),
	.datab(av_readdata_pre_21),
	.datac(gnd),
	.datad(\wb_dmem_read_data[7]~17_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data[5]~3_combout ),
	.cout());
defparam \wb_dmem_read_data[5]~3 .lut_mask = 16'hCCAA;
defparam \wb_dmem_read_data[5]~3 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[5] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data[5]~3_combout ),
	.asdata(av_readdata_pre_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\wb_dmem_read_data[7]~19_combout ),
	.sload(\wb_dmem_read_data[7]~21_combout ),
	.ena(vcc),
	.q(\wb_dmem_read_data[5]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[5] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[5] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[5]~46 (
	.dataa(\wb_npc[5]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[5]~45_combout ),
	.datad(\wb_dmem_read_data[5]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[5]~46_combout ),
	.cout());
defparam \_T_3543__T_3854_data[5]~46 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[5]~46 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a27 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[5]~46_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a27_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_a_first_bit_number = 27;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_b_first_bit_number = 27;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a27 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~22 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a27~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~22_combout ),
	.cout());
defparam \ex_rs_0~22 .lut_mask = 16'h0080;
defparam \ex_rs_0~22 .sum_lutc_input = "datac";

dffeas \ex_rs_0[5] (
	.clk(clk_clk),
	.d(\ex_rs_0~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[5]~q ),
	.prn(vcc));
defparam \ex_rs_0[5] .is_wysiwyg = "true";
defparam \ex_rs_0[5] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[5]~91 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(\ex_rs_0[5]~q ),
	.datac(\wb_alu_out[5]~q ),
	.datad(\ex_reg_rs1_bypass[2]~7_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[5]~91_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[5]~91 .lut_mask = 16'hAAD8;
defparam \ex_reg_rs1_bypass[5]~91 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[5]~92 (
	.dataa(av_readdata_pre_5),
	.datab(\wb_csr_data[5]~q ),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\ex_reg_rs1_bypass[5]~91_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[5]~92_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[5]~92 .lut_mask = 16'hCFA0;
defparam \ex_reg_rs1_bypass[5]~92 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[5]~93 (
	.dataa(\ex_reg_rs1_bypass[0]~4_combout ),
	.datab(\ex_reg_rs1_bypass[5]~90_combout ),
	.datac(\ex_reg_rs1_bypass[5]~92_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[5]~93_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[5]~93 .lut_mask = 16'hECEC;
defparam \ex_reg_rs1_bypass[5]~93 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[5]~108 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[5]~q ),
	.datad(\ex_reg_rs1_bypass[5]~93_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[5]~108_combout ),
	.cout());
defparam \alu_io_op1[5]~108 .lut_mask = 16'h6240;
defparam \alu_io_op1[5]~108 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[5]~43 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_ctrl_imm_type.101~q ),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\alu_io_op2[5]~43_combout ),
	.cout());
defparam \alu_io_op2[5]~43 .lut_mask = 16'h888B;
defparam \alu_io_op2[5]~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_csr_addr~9 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[25]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_csr_addr~9_combout ),
	.cout());
defparam \ex_csr_addr~9 .lut_mask = 16'h8080;
defparam \ex_csr_addr~9 .sum_lutc_input = "datac";

dffeas \ex_csr_addr[5] (
	.clk(clk_clk),
	.d(\ex_csr_addr~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_addr[5]~q ),
	.prn(vcc));
defparam \ex_csr_addr[5] .is_wysiwyg = "true";
defparam \ex_csr_addr[5] .power_up = "low";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a27 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[5]~46_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a27_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_a_first_bit_number = 27;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_b_first_bit_number = 27;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a27 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~23 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a27~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~23_combout ),
	.cout());
defparam \ex_rs_1~23 .lut_mask = 16'h8888;
defparam \ex_rs_1~23 .sum_lutc_input = "datac";

dffeas \ex_rs_1[5] (
	.clk(clk_clk),
	.d(\ex_rs_1~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[5]~q ),
	.prn(vcc));
defparam \ex_rs_1[5] .is_wysiwyg = "true";
defparam \ex_rs_1[5] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[5]~83 (
	.dataa(\ex_reg_rs2_bypass[7]~5_combout ),
	.datab(\ex_rs_1[5]~q ),
	.datac(\ex_reg_rs2_bypass[7]~4_combout ),
	.datad(\wb_alu_out[5]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[5]~83_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[5]~83 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[5]~83 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[5]~84 (
	.dataa(av_readdata_pre_5),
	.datab(\ex_reg_rs2_bypass[7]~5_combout ),
	.datac(\ex_reg_rs2_bypass[5]~83_combout ),
	.datad(\wb_csr_data[5]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[5]~84_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[5]~84 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[5]~84 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[5]~85 (
	.dataa(\mem_alu_out[5]~q ),
	.datab(\ex_reg_rs2_bypass[5]~84_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[5]~85_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[5]~85 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[5]~85 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[5]~67 (
	.dataa(\_T_3681~3_combout ),
	.datab(\mem_csr_data[5]~q ),
	.datac(\ex_reg_rs2_bypass[5]~85_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\alu_io_op2[5]~67_combout ),
	.cout());
defparam \alu_io_op2[5]~67 .lut_mask = 16'hF8F8;
defparam \alu_io_op2[5]~67 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[5]~68 (
	.dataa(\alu_io_op2[5]~43_combout ),
	.datab(\ex_csr_addr[5]~q ),
	.datac(\ex_ctrl_alu_op2.10~q ),
	.datad(\alu_io_op2[5]~67_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[5]~68_combout ),
	.cout());
defparam \alu_io_op2[5]~68 .lut_mask = 16'hA808;
defparam \alu_io_op2[5]~68 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~141 (
	.dataa(\mem_alu_out[26]~2_combout ),
	.datab(\alu|LessThan0~0_combout ),
	.datac(\alu_io_op2[5]~68_combout ),
	.datad(\alu_io_op1[5]~108_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~141_combout ),
	.cout());
defparam \mem_alu_out~141 .lut_mask = 16'h7DD4;
defparam \mem_alu_out~141 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~142 (
	.dataa(\mem_alu_out[26]~2_combout ),
	.datab(\mem_alu_out~141_combout ),
	.datac(\alu|LessThan0~0_combout ),
	.datad(\alu|ShiftRight0~253_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~142_combout ),
	.cout());
defparam \mem_alu_out~142 .lut_mask = 16'hCC8C;
defparam \mem_alu_out~142 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~88 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[5]~68_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~142_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~88_combout ),
	.cout());
defparam \mem_alu_out~88 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~88 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~89 (
	.dataa(\alu_io_op1[5]~108_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~88_combout ),
	.datad(\alu|ShiftRight0~233_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~89_combout ),
	.cout());
defparam \mem_alu_out~89 .lut_mask = 16'hF838;
defparam \mem_alu_out~89 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~90 (
	.dataa(\mem_alu_out~89_combout ),
	.datab(\alu|_T_3[5]~10_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~90_combout ),
	.cout());
defparam \mem_alu_out~90 .lut_mask = 16'h00AC;
defparam \mem_alu_out~90 .sum_lutc_input = "datac";

dffeas \mem_alu_out[5] (
	.clk(clk_clk),
	.d(\mem_alu_out~90_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[5]~q ),
	.prn(vcc));
defparam \mem_alu_out[5] .is_wysiwyg = "true";
defparam \mem_alu_out[5] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~3 (
	.dataa(\ex_pc[5]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~3_combout ),
	.cout());
defparam \mem_pc~3 .lut_mask = 16'h8888;
defparam \mem_pc~3 .sum_lutc_input = "datac";

dffeas \mem_pc[5] (
	.clk(clk_clk),
	.d(\mem_pc~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[5]~q ),
	.prn(vcc));
defparam \mem_pc[5] .is_wysiwyg = "true";
defparam \mem_pc[5] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~20 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_csr_addr[5]~q ),
	.datac(\ex_ctrl_imm_type.101~q ),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\mem_imm~20_combout ),
	.cout());
defparam \mem_imm~20 .lut_mask = 16'h0008;
defparam \mem_imm~20 .sum_lutc_input = "datac";

dffeas \mem_imm[5] (
	.clk(clk_clk),
	.d(\mem_imm~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[5]~q ),
	.prn(vcc));
defparam \mem_imm[5] .is_wysiwyg = "true";
defparam \mem_imm[5] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[5]~10 (
	.dataa(\mem_pc[5]~q ),
	.datab(\mem_imm[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[4]~9 ),
	.combout(\_T_3862[5]~10_combout ),
	.cout(\_T_3862[5]~11 ));
defparam \_T_3862[5]~10 .lut_mask = 16'h9617;
defparam \_T_3862[5]~10 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~19 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[5]~10_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[5]~6_combout ),
	.cin(gnd),
	.combout(\pc_cntr~19_combout ),
	.cout());
defparam \pc_cntr~19 .lut_mask = 16'h5E0E;
defparam \pc_cntr~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~20 (
	.dataa(\mem_alu_out[5]~q ),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~19_combout ),
	.datad(\csr|mepc[5]~q ),
	.cin(gnd),
	.combout(\pc_cntr~20_combout ),
	.cout());
defparam \pc_cntr~20 .lut_mask = 16'hF838;
defparam \pc_cntr~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~21 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~20_combout ),
	.datac(\csr|mtvec[5]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~21_combout ),
	.cout());
defparam \pc_cntr~21 .lut_mask = 16'h88A0;
defparam \pc_cntr~21 .sum_lutc_input = "datac";

dffeas \pc_cntr[5] (
	.clk(clk_clk),
	.d(\pc_cntr~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[5]~q ),
	.prn(vcc));
defparam \pc_cntr[5] .is_wysiwyg = "true";
defparam \pc_cntr[5] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~4 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~4_combout ),
	.cout());
defparam \id_pc~4 .lut_mask = 16'h8080;
defparam \id_pc~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~2 (
	.dataa(id_pc_6),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~2_combout ),
	.cout());
defparam \ex_pc~2 .lut_mask = 16'h8080;
defparam \ex_pc~2 .sum_lutc_input = "datac";

dffeas \ex_pc[6] (
	.clk(clk_clk),
	.d(\ex_pc~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[6]~q ),
	.prn(vcc));
defparam \ex_pc[6] .is_wysiwyg = "true";
defparam \ex_pc[6] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~4 (
	.dataa(\ex_pc[6]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~4_combout ),
	.cout());
defparam \mem_pc~4 .lut_mask = 16'h8888;
defparam \mem_pc~4 .sum_lutc_input = "datac";

dffeas \mem_pc[6] (
	.clk(clk_clk),
	.d(\mem_pc~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[6]~q ),
	.prn(vcc));
defparam \mem_pc[6] .is_wysiwyg = "true";
defparam \mem_pc[6] .power_up = "low";

cyclone10lp_lcell_comb \ex_csr_addr~10 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[26]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_csr_addr~10_combout ),
	.cout());
defparam \ex_csr_addr~10 .lut_mask = 16'h8080;
defparam \ex_csr_addr~10 .sum_lutc_input = "datac";

dffeas \ex_csr_addr[6] (
	.clk(clk_clk),
	.d(\ex_csr_addr~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_addr[6]~q ),
	.prn(vcc));
defparam \ex_csr_addr[6] .is_wysiwyg = "true";
defparam \ex_csr_addr[6] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~21 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_csr_addr[6]~q ),
	.datac(\ex_ctrl_imm_type.101~q ),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\mem_imm~21_combout ),
	.cout());
defparam \mem_imm~21 .lut_mask = 16'h0008;
defparam \mem_imm~21 .sum_lutc_input = "datac";

dffeas \mem_imm[6] (
	.clk(clk_clk),
	.d(\mem_imm~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[6]~q ),
	.prn(vcc));
defparam \mem_imm[6] .is_wysiwyg = "true";
defparam \mem_imm[6] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[6]~12 (
	.dataa(\mem_pc[6]~q ),
	.datab(\mem_imm[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[5]~11 ),
	.combout(\_T_3862[6]~12_combout ),
	.cout(\_T_3862[6]~13 ));
defparam \_T_3862[6]~12 .lut_mask = 16'h698E;
defparam \_T_3862[6]~12 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \mem_csr_data~29 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[6]~173_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~29_combout ),
	.cout());
defparam \mem_csr_data~29 .lut_mask = 16'h8888;
defparam \mem_csr_data~29 .sum_lutc_input = "datac";

dffeas \mem_csr_data[6] (
	.clk(clk_clk),
	.d(\mem_csr_data~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[6]~q ),
	.prn(vcc));
defparam \mem_csr_data[6] .is_wysiwyg = "true";
defparam \mem_csr_data[6] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~22 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~22_combout ),
	.cout());
defparam \wb_csr_data~22 .lut_mask = 16'h8888;
defparam \wb_csr_data~22 .sum_lutc_input = "datac";

dffeas \wb_csr_data[6] (
	.clk(clk_clk),
	.d(\wb_csr_data~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[6]~q ),
	.prn(vcc));
defparam \wb_csr_data[6] .is_wysiwyg = "true";
defparam \wb_csr_data[6] .power_up = "low";

cyclone10lp_lcell_comb \npc[6]~8 (
	.dataa(\pc_cntr[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[5]~7 ),
	.combout(\npc[6]~8_combout ),
	.cout(\npc[6]~9 ));
defparam \npc[6]~8 .lut_mask = 16'hA50A;
defparam \npc[6]~8 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~22 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[6]~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~22_combout ),
	.cout());
defparam \id_npc~22 .lut_mask = 16'h8080;
defparam \id_npc~22 .sum_lutc_input = "datac";

dffeas \id_npc[6] (
	.clk(clk_clk),
	.d(\id_npc~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[6]~q ),
	.prn(vcc));
defparam \id_npc[6] .is_wysiwyg = "true";
defparam \id_npc[6] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~22 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[6]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~22_combout ),
	.cout());
defparam \ex_npc~22 .lut_mask = 16'h8080;
defparam \ex_npc~22 .sum_lutc_input = "datac";

dffeas \ex_npc[6] (
	.clk(clk_clk),
	.d(\ex_npc~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[6]~q ),
	.prn(vcc));
defparam \ex_npc[6] .is_wysiwyg = "true";
defparam \ex_npc[6] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~20 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~20_combout ),
	.cout());
defparam \mem_npc~20 .lut_mask = 16'h8888;
defparam \mem_npc~20 .sum_lutc_input = "datac";

dffeas \mem_npc[6] (
	.clk(clk_clk),
	.d(\mem_npc~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[6]~q ),
	.prn(vcc));
defparam \mem_npc[6] .is_wysiwyg = "true";
defparam \mem_npc[6] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~20 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~20_combout ),
	.cout());
defparam \wb_npc~20 .lut_mask = 16'h8888;
defparam \wb_npc~20 .sum_lutc_input = "datac";

dffeas \wb_npc[6] (
	.clk(clk_clk),
	.d(\wb_npc~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[6]~q ),
	.prn(vcc));
defparam \wb_npc[6] .is_wysiwyg = "true";
defparam \wb_npc[6] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~22 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~22_combout ),
	.cout());
defparam \wb_alu_out~22 .lut_mask = 16'h8888;
defparam \wb_alu_out~22 .sum_lutc_input = "datac";

dffeas \wb_alu_out[6] (
	.clk(clk_clk),
	.d(\wb_alu_out~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[6]~q ),
	.prn(vcc));
defparam \wb_alu_out[6] .is_wysiwyg = "true";
defparam \wb_alu_out[6] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[6]~47 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[6]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[6]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[6]~47_combout ),
	.cout());
defparam \_T_3543__T_3854_data[6]~47 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[6]~47 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~68 (
	.dataa(av_readdata_pre_30),
	.datab(av_readdata_pre_14),
	.datac(gnd),
	.datad(mem_alu_out_1),
	.cin(gnd),
	.combout(\wb_dmem_read_data~68_combout ),
	.cout());
defparam \wb_dmem_read_data~68 .lut_mask = 16'hAACC;
defparam \wb_dmem_read_data~68 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[6]~2 (
	.dataa(\wb_dmem_read_data~68_combout ),
	.datab(av_readdata_pre_22),
	.datac(gnd),
	.datad(\wb_dmem_read_data[7]~17_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data[6]~2_combout ),
	.cout());
defparam \wb_dmem_read_data[6]~2 .lut_mask = 16'hCCAA;
defparam \wb_dmem_read_data[6]~2 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[6] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data[6]~2_combout ),
	.asdata(av_readdata_pre_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\wb_dmem_read_data[7]~19_combout ),
	.sload(\wb_dmem_read_data[7]~21_combout ),
	.ena(vcc),
	.q(\wb_dmem_read_data[6]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[6] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[6] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[6]~48 (
	.dataa(\wb_csr_data[6]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[6]~47_combout ),
	.datad(\wb_dmem_read_data[6]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[6]~48_combout ),
	.cout());
defparam \_T_3543__T_3854_data[6]~48 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[6]~48 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a26 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[6]~48_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a26_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_a_first_bit_number = 26;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_b_first_bit_number = 26;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a26 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~24 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a26~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~24_combout ),
	.cout());
defparam \ex_rs_1~24 .lut_mask = 16'h8888;
defparam \ex_rs_1~24 .sum_lutc_input = "datac";

dffeas \ex_rs_1[6] (
	.clk(clk_clk),
	.d(\ex_rs_1~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[6]~q ),
	.prn(vcc));
defparam \ex_rs_1[6] .is_wysiwyg = "true";
defparam \ex_rs_1[6] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[6]~86 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_6),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[6]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[6]~86_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[6]~86 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[6]~86 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[6]~87 (
	.dataa(\ex_rs_1[6]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[6]~86_combout ),
	.datad(\wb_csr_data[6]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[6]~87_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[6]~87 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[6]~87 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[6]~88 (
	.dataa(\mem_alu_out[6]~q ),
	.datab(\ex_reg_rs2_bypass[6]~87_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[6]~88_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[6]~88 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[6]~88 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[6]~69 (
	.dataa(\_T_3681~3_combout ),
	.datab(\mem_csr_data[6]~q ),
	.datac(\ex_reg_rs2_bypass[6]~88_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\alu_io_op2[6]~69_combout ),
	.cout());
defparam \alu_io_op2[6]~69 .lut_mask = 16'hF8F8;
defparam \alu_io_op2[6]~69 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[6]~70 (
	.dataa(\alu_io_op2[5]~43_combout ),
	.datab(\ex_csr_addr[6]~q ),
	.datac(\ex_ctrl_alu_op2.10~q ),
	.datad(\alu_io_op2[6]~69_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[6]~70_combout ),
	.cout());
defparam \alu_io_op2[6]~70 .lut_mask = 16'hA808;
defparam \alu_io_op2[6]~70 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[6]~98 (
	.dataa(\ex_reg_rs1_bypass[0]~20_combout ),
	.datab(\mem_alu_out[6]~q ),
	.datac(\_T_3634~2_combout ),
	.datad(\mem_csr_data[6]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[6]~98_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[6]~98 .lut_mask = 16'hF888;
defparam \ex_reg_rs1_bypass[6]~98 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a26 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[6]~48_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a26_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_a_first_bit_number = 26;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_b_first_bit_number = 26;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a26 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~24 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a26~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~24_combout ),
	.cout());
defparam \ex_rs_0~24 .lut_mask = 16'h0080;
defparam \ex_rs_0~24 .sum_lutc_input = "datac";

dffeas \ex_rs_0[6] (
	.clk(clk_clk),
	.d(\ex_rs_0~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[6]~q ),
	.prn(vcc));
defparam \ex_rs_0[6] .is_wysiwyg = "true";
defparam \ex_rs_0[6] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[6]~99 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(av_readdata_pre_6),
	.datac(\wb_alu_out[6]~q ),
	.datad(\ex_reg_rs1_bypass[2]~138_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[6]~99_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[6]~99 .lut_mask = 16'hAAD8;
defparam \ex_reg_rs1_bypass[6]~99 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[6]~100 (
	.dataa(\ex_rs_0[6]~q ),
	.datab(\wb_csr_data[6]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\ex_reg_rs1_bypass[6]~99_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[6]~100_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[6]~100 .lut_mask = 16'hCFA0;
defparam \ex_reg_rs1_bypass[6]~100 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[6]~101 (
	.dataa(\ex_reg_rs1_bypass[0]~4_combout ),
	.datab(\ex_reg_rs1_bypass[6]~98_combout ),
	.datac(\ex_reg_rs1_bypass[6]~100_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[6]~101_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[6]~101 .lut_mask = 16'hECEC;
defparam \ex_reg_rs1_bypass[6]~101 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[6]~110 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[6]~q ),
	.datad(\ex_reg_rs1_bypass[6]~101_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[6]~110_combout ),
	.cout());
defparam \alu_io_op1[6]~110 .lut_mask = 16'h6240;
defparam \alu_io_op1[6]~110 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~139 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\alu_io_op2[6]~70_combout ),
	.datad(\alu_io_op1[6]~110_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~139_combout ),
	.cout());
defparam \mem_alu_out~139 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~139 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~140 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~139_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~254_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~140_combout ),
	.cout());
defparam \mem_alu_out~140 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~140 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~91 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[6]~110_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~140_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~91_combout ),
	.cout());
defparam \mem_alu_out~91 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~91 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~92 (
	.dataa(\alu_io_op2[6]~70_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~91_combout ),
	.datad(\alu|ShiftRight0~236_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~92_combout ),
	.cout());
defparam \mem_alu_out~92 .lut_mask = 16'hF838;
defparam \mem_alu_out~92 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~93 (
	.dataa(\mem_alu_out~92_combout ),
	.datab(\alu|_T_3[6]~12_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~93_combout ),
	.cout());
defparam \mem_alu_out~93 .lut_mask = 16'h00AC;
defparam \mem_alu_out~93 .sum_lutc_input = "datac";

dffeas \mem_alu_out[6] (
	.clk(clk_clk),
	.d(\mem_alu_out~93_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[6]~q ),
	.prn(vcc));
defparam \mem_alu_out[6] .is_wysiwyg = "true";
defparam \mem_alu_out[6] .power_up = "low";

cyclone10lp_lcell_comb \pc_cntr~22 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(\mem_alu_out[6]~q ),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[6]~8_combout ),
	.cin(gnd),
	.combout(\pc_cntr~22_combout ),
	.cout());
defparam \pc_cntr~22 .lut_mask = 16'hDAD0;
defparam \pc_cntr~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~23 (
	.dataa(\_T_3862[6]~12_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~22_combout ),
	.datad(\csr|mepc[6]~q ),
	.cin(gnd),
	.combout(\pc_cntr~23_combout ),
	.cout());
defparam \pc_cntr~23 .lut_mask = 16'hF2C2;
defparam \pc_cntr~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~24 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~23_combout ),
	.datac(\csr|mtvec[6]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~24_combout ),
	.cout());
defparam \pc_cntr~24 .lut_mask = 16'h88A0;
defparam \pc_cntr~24 .sum_lutc_input = "datac";

dffeas \pc_cntr[6] (
	.clk(clk_clk),
	.d(\pc_cntr~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[6]~q ),
	.prn(vcc));
defparam \pc_cntr[6] .is_wysiwyg = "true";
defparam \pc_cntr[6] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~5 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[6]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~5_combout ),
	.cout());
defparam \id_pc~5 .lut_mask = 16'h8080;
defparam \id_pc~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~3 (
	.dataa(id_pc_7),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~3_combout ),
	.cout());
defparam \ex_pc~3 .lut_mask = 16'h8080;
defparam \ex_pc~3 .sum_lutc_input = "datac";

dffeas \ex_pc[7] (
	.clk(clk_clk),
	.d(\ex_pc~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[7]~q ),
	.prn(vcc));
defparam \ex_pc[7] .is_wysiwyg = "true";
defparam \ex_pc[7] .power_up = "low";

cyclone10lp_lcell_comb \mem_csr_data~30 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[7]~181_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~30_combout ),
	.cout());
defparam \mem_csr_data~30 .lut_mask = 16'h8888;
defparam \mem_csr_data~30 .sum_lutc_input = "datac";

dffeas \mem_csr_data[7] (
	.clk(clk_clk),
	.d(\mem_csr_data~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[7]~q ),
	.prn(vcc));
defparam \mem_csr_data[7] .is_wysiwyg = "true";
defparam \mem_csr_data[7] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[7]~102 (
	.dataa(\ex_reg_rs1_bypass[0]~20_combout ),
	.datab(\mem_alu_out[7]~q ),
	.datac(\_T_3634~2_combout ),
	.datad(\mem_csr_data[7]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[7]~102_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[7]~102 .lut_mask = 16'hF888;
defparam \ex_reg_rs1_bypass[7]~102 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_csr_data~23 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~23_combout ),
	.cout());
defparam \wb_csr_data~23 .lut_mask = 16'h8888;
defparam \wb_csr_data~23 .sum_lutc_input = "datac";

dffeas \wb_csr_data[7] (
	.clk(clk_clk),
	.d(\wb_csr_data~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[7]~q ),
	.prn(vcc));
defparam \wb_csr_data[7] .is_wysiwyg = "true";
defparam \wb_csr_data[7] .power_up = "low";

cyclone10lp_lcell_comb \npc[7]~10 (
	.dataa(\pc_cntr[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[6]~9 ),
	.combout(\npc[7]~10_combout ),
	.cout(\npc[7]~11 ));
defparam \npc[7]~10 .lut_mask = 16'h5A5F;
defparam \npc[7]~10 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~23 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[7]~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~23_combout ),
	.cout());
defparam \id_npc~23 .lut_mask = 16'h8080;
defparam \id_npc~23 .sum_lutc_input = "datac";

dffeas \id_npc[7] (
	.clk(clk_clk),
	.d(\id_npc~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[7]~q ),
	.prn(vcc));
defparam \id_npc[7] .is_wysiwyg = "true";
defparam \id_npc[7] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~23 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~23_combout ),
	.cout());
defparam \ex_npc~23 .lut_mask = 16'h8080;
defparam \ex_npc~23 .sum_lutc_input = "datac";

dffeas \ex_npc[7] (
	.clk(clk_clk),
	.d(\ex_npc~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[7]~q ),
	.prn(vcc));
defparam \ex_npc[7] .is_wysiwyg = "true";
defparam \ex_npc[7] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~21 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~21_combout ),
	.cout());
defparam \mem_npc~21 .lut_mask = 16'h8888;
defparam \mem_npc~21 .sum_lutc_input = "datac";

dffeas \mem_npc[7] (
	.clk(clk_clk),
	.d(\mem_npc~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[7]~q ),
	.prn(vcc));
defparam \mem_npc[7] .is_wysiwyg = "true";
defparam \mem_npc[7] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~21 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~21_combout ),
	.cout());
defparam \wb_npc~21 .lut_mask = 16'h8888;
defparam \wb_npc~21 .sum_lutc_input = "datac";

dffeas \wb_npc[7] (
	.clk(clk_clk),
	.d(\wb_npc~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[7]~q ),
	.prn(vcc));
defparam \wb_npc[7] .is_wysiwyg = "true";
defparam \wb_npc[7] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~23 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~23_combout ),
	.cout());
defparam \wb_alu_out~23 .lut_mask = 16'h8888;
defparam \wb_alu_out~23 .sum_lutc_input = "datac";

dffeas \wb_alu_out[7] (
	.clk(clk_clk),
	.d(\wb_alu_out~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[7]~q ),
	.prn(vcc));
defparam \wb_alu_out[7] .is_wysiwyg = "true";
defparam \wb_alu_out[7] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[7]~49 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[7]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[7]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[7]~49_combout ),
	.cout());
defparam \_T_3543__T_3854_data[7]~49 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[7]~49 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~28 (
	.dataa(av_readdata_pre_31),
	.datab(av_readdata_pre_15),
	.datac(gnd),
	.datad(mem_alu_out_1),
	.cin(gnd),
	.combout(\wb_dmem_read_data~28_combout ),
	.cout());
defparam \wb_dmem_read_data~28 .lut_mask = 16'hAACC;
defparam \wb_dmem_read_data~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[7]~1 (
	.dataa(\wb_dmem_read_data~28_combout ),
	.datab(av_readdata_pre_23),
	.datac(gnd),
	.datad(\wb_dmem_read_data[7]~17_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data[7]~1_combout ),
	.cout());
defparam \wb_dmem_read_data[7]~1 .lut_mask = 16'hCCAA;
defparam \wb_dmem_read_data[7]~1 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[7] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data[7]~1_combout ),
	.asdata(av_readdata_pre_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\wb_dmem_read_data[7]~19_combout ),
	.sload(\wb_dmem_read_data[7]~21_combout ),
	.ena(vcc),
	.q(\wb_dmem_read_data[7]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[7] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[7] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[7]~50 (
	.dataa(\wb_npc[7]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[7]~49_combout ),
	.datad(\wb_dmem_read_data[7]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[7]~50_combout ),
	.cout());
defparam \_T_3543__T_3854_data[7]~50 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[7]~50 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a25 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[7]~50_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a25_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_a_first_bit_number = 25;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_b_first_bit_number = 25;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a25 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~25 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a25~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~25_combout ),
	.cout());
defparam \ex_rs_0~25 .lut_mask = 16'h0080;
defparam \ex_rs_0~25 .sum_lutc_input = "datac";

dffeas \ex_rs_0[7] (
	.clk(clk_clk),
	.d(\ex_rs_0~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[7]~q ),
	.prn(vcc));
defparam \ex_rs_0[7] .is_wysiwyg = "true";
defparam \ex_rs_0[7] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[7]~103 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(\ex_rs_0[7]~q ),
	.datac(\wb_alu_out[7]~q ),
	.datad(\ex_reg_rs1_bypass[2]~7_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[7]~103_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[7]~103 .lut_mask = 16'hAAD8;
defparam \ex_reg_rs1_bypass[7]~103 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[7]~104 (
	.dataa(av_readdata_pre_7),
	.datab(\wb_csr_data[7]~q ),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\ex_reg_rs1_bypass[7]~103_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[7]~104_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[7]~104 .lut_mask = 16'hCFA0;
defparam \ex_reg_rs1_bypass[7]~104 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[7]~105 (
	.dataa(\ex_reg_rs1_bypass[0]~4_combout ),
	.datab(\ex_reg_rs1_bypass[7]~102_combout ),
	.datac(\ex_reg_rs1_bypass[7]~104_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[7]~105_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[7]~105 .lut_mask = 16'hECEC;
defparam \ex_reg_rs1_bypass[7]~105 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[7]~111 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[7]~q ),
	.datad(\ex_reg_rs1_bypass[7]~105_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[7]~111_combout ),
	.cout());
defparam \alu_io_op1[7]~111 .lut_mask = 16'h6240;
defparam \alu_io_op1[7]~111 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_csr_addr~11 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[27]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_csr_addr~11_combout ),
	.cout());
defparam \ex_csr_addr~11 .lut_mask = 16'h8080;
defparam \ex_csr_addr~11 .sum_lutc_input = "datac";

dffeas \ex_csr_addr[7] (
	.clk(clk_clk),
	.d(\ex_csr_addr~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_addr[7]~q ),
	.prn(vcc));
defparam \ex_csr_addr[7] .is_wysiwyg = "true";
defparam \ex_csr_addr[7] .power_up = "low";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a25 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[7]~50_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a25_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_a_first_bit_number = 25;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_b_first_bit_number = 25;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a25 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~25 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a25~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~25_combout ),
	.cout());
defparam \ex_rs_1~25 .lut_mask = 16'h8888;
defparam \ex_rs_1~25 .sum_lutc_input = "datac";

dffeas \ex_rs_1[7] (
	.clk(clk_clk),
	.d(\ex_rs_1~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[7]~q ),
	.prn(vcc));
defparam \ex_rs_1[7] .is_wysiwyg = "true";
defparam \ex_rs_1[7] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[7]~89 (
	.dataa(\ex_reg_rs2_bypass[7]~5_combout ),
	.datab(\ex_rs_1[7]~q ),
	.datac(\ex_reg_rs2_bypass[7]~4_combout ),
	.datad(\wb_alu_out[7]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[7]~89_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[7]~89 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[7]~89 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[7]~90 (
	.dataa(av_readdata_pre_7),
	.datab(\ex_reg_rs2_bypass[7]~5_combout ),
	.datac(\ex_reg_rs2_bypass[7]~89_combout ),
	.datad(\wb_csr_data[7]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[7]~90_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[7]~90 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[7]~90 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[7]~91 (
	.dataa(\mem_alu_out[7]~q ),
	.datab(\ex_reg_rs2_bypass[7]~90_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[7]~91_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[7]~91 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[7]~91 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[7]~71 (
	.dataa(\_T_3681~3_combout ),
	.datab(\mem_csr_data[7]~q ),
	.datac(\ex_reg_rs2_bypass[7]~91_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\alu_io_op2[7]~71_combout ),
	.cout());
defparam \alu_io_op2[7]~71 .lut_mask = 16'hF8F8;
defparam \alu_io_op2[7]~71 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[7]~72 (
	.dataa(\alu_io_op2[5]~43_combout ),
	.datab(\ex_csr_addr[7]~q ),
	.datac(\ex_ctrl_alu_op2.10~q ),
	.datad(\alu_io_op2[7]~71_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[7]~72_combout ),
	.cout());
defparam \alu_io_op2[7]~72 .lut_mask = 16'hA808;
defparam \alu_io_op2[7]~72 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~94 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\alu|_T_123[7]~combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~256_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~94_combout ),
	.cout());
defparam \mem_alu_out~94 .lut_mask = 16'hDAD0;
defparam \mem_alu_out~94 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~95 (
	.dataa(\alu_io_op1[7]~111_combout ),
	.datab(\alu_io_op2[7]~72_combout ),
	.datac(\mem_alu_out~94_combout ),
	.datad(\alu|LessThan0~0_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~95_combout ),
	.cout());
defparam \mem_alu_out~95 .lut_mask = 16'hF08E;
defparam \mem_alu_out~95 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~96 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[7]~72_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~95_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~96_combout ),
	.cout());
defparam \mem_alu_out~96 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~96 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~97 (
	.dataa(\alu_io_op1[7]~111_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~96_combout ),
	.datad(\alu|ShiftRight0~240_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~97_combout ),
	.cout());
defparam \mem_alu_out~97 .lut_mask = 16'hF838;
defparam \mem_alu_out~97 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~98 (
	.dataa(\mem_alu_out~97_combout ),
	.datab(\alu|_T_3[7]~14_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~98_combout ),
	.cout());
defparam \mem_alu_out~98 .lut_mask = 16'h00AC;
defparam \mem_alu_out~98 .sum_lutc_input = "datac";

dffeas \mem_alu_out[7] (
	.clk(clk_clk),
	.d(\mem_alu_out~98_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[7]~q ),
	.prn(vcc));
defparam \mem_alu_out[7] .is_wysiwyg = "true";
defparam \mem_alu_out[7] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~5 (
	.dataa(\ex_pc[7]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~5_combout ),
	.cout());
defparam \mem_pc~5 .lut_mask = 16'h8888;
defparam \mem_pc~5 .sum_lutc_input = "datac";

dffeas \mem_pc[7] (
	.clk(clk_clk),
	.d(\mem_pc~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[7]~q ),
	.prn(vcc));
defparam \mem_pc[7] .is_wysiwyg = "true";
defparam \mem_pc[7] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~22 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_csr_addr[7]~q ),
	.datac(\ex_ctrl_imm_type.101~q ),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\mem_imm~22_combout ),
	.cout());
defparam \mem_imm~22 .lut_mask = 16'h0008;
defparam \mem_imm~22 .sum_lutc_input = "datac";

dffeas \mem_imm[7] (
	.clk(clk_clk),
	.d(\mem_imm~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[7]~q ),
	.prn(vcc));
defparam \mem_imm[7] .is_wysiwyg = "true";
defparam \mem_imm[7] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[7]~14 (
	.dataa(\mem_pc[7]~q ),
	.datab(\mem_imm[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[6]~13 ),
	.combout(\_T_3862[7]~14_combout ),
	.cout(\_T_3862[7]~15 ));
defparam \_T_3862[7]~14 .lut_mask = 16'h9617;
defparam \_T_3862[7]~14 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~25 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[7]~14_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[7]~10_combout ),
	.cin(gnd),
	.combout(\pc_cntr~25_combout ),
	.cout());
defparam \pc_cntr~25 .lut_mask = 16'h5E0E;
defparam \pc_cntr~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~26 (
	.dataa(\mem_alu_out[7]~q ),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~25_combout ),
	.datad(\csr|mepc[7]~q ),
	.cin(gnd),
	.combout(\pc_cntr~26_combout ),
	.cout());
defparam \pc_cntr~26 .lut_mask = 16'hF838;
defparam \pc_cntr~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~27 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~26_combout ),
	.datac(\csr|mtvec[7]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~27_combout ),
	.cout());
defparam \pc_cntr~27 .lut_mask = 16'h88A0;
defparam \pc_cntr~27 .sum_lutc_input = "datac";

dffeas \pc_cntr[7] (
	.clk(clk_clk),
	.d(\pc_cntr~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[7]~q ),
	.prn(vcc));
defparam \pc_cntr[7] .is_wysiwyg = "true";
defparam \pc_cntr[7] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~6 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~6_combout ),
	.cout());
defparam \id_pc~6 .lut_mask = 16'h8080;
defparam \id_pc~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~6 (
	.dataa(id_pc_8),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~6_combout ),
	.cout());
defparam \ex_pc~6 .lut_mask = 16'h8080;
defparam \ex_pc~6 .sum_lutc_input = "datac";

dffeas \ex_pc[8] (
	.clk(clk_clk),
	.d(\ex_pc~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[8]~q ),
	.prn(vcc));
defparam \ex_pc[8] .is_wysiwyg = "true";
defparam \ex_pc[8] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~6 (
	.dataa(\ex_pc[8]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~6_combout ),
	.cout());
defparam \mem_pc~6 .lut_mask = 16'h8888;
defparam \mem_pc~6 .sum_lutc_input = "datac";

dffeas \mem_pc[8] (
	.clk(clk_clk),
	.d(\mem_pc~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[8]~q ),
	.prn(vcc));
defparam \mem_pc[8] .is_wysiwyg = "true";
defparam \mem_pc[8] .power_up = "low";

cyclone10lp_lcell_comb \ex_csr_addr~5 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[28]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_csr_addr~5_combout ),
	.cout());
defparam \ex_csr_addr~5 .lut_mask = 16'h8080;
defparam \ex_csr_addr~5 .sum_lutc_input = "datac";

dffeas \ex_csr_addr[8] (
	.clk(clk_clk),
	.d(\ex_csr_addr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_addr[8]~q ),
	.prn(vcc));
defparam \ex_csr_addr[8] .is_wysiwyg = "true";
defparam \ex_csr_addr[8] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~23 (
	.dataa(\ex_csr_addr[8]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(\ex_ctrl_imm_type.101~q ),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\mem_imm~23_combout ),
	.cout());
defparam \mem_imm~23 .lut_mask = 16'h0008;
defparam \mem_imm~23 .sum_lutc_input = "datac";

dffeas \mem_imm[8] (
	.clk(clk_clk),
	.d(\mem_imm~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[8]~q ),
	.prn(vcc));
defparam \mem_imm[8] .is_wysiwyg = "true";
defparam \mem_imm[8] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[8]~16 (
	.dataa(\mem_pc[8]~q ),
	.datab(\mem_imm[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[7]~15 ),
	.combout(\_T_3862[8]~16_combout ),
	.cout(\_T_3862[8]~17 ));
defparam \_T_3862[8]~16 .lut_mask = 16'h698E;
defparam \_T_3862[8]~16 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \mem_csr_data~13 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[8]~59_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~13_combout ),
	.cout());
defparam \mem_csr_data~13 .lut_mask = 16'h8888;
defparam \mem_csr_data~13 .sum_lutc_input = "datac";

dffeas \mem_csr_data[8] (
	.clk(clk_clk),
	.d(\mem_csr_data~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[8]~q ),
	.prn(vcc));
defparam \mem_csr_data[8] .is_wysiwyg = "true";
defparam \mem_csr_data[8] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~6 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~6_combout ),
	.cout());
defparam \wb_csr_data~6 .lut_mask = 16'h8888;
defparam \wb_csr_data~6 .sum_lutc_input = "datac";

dffeas \wb_csr_data[8] (
	.clk(clk_clk),
	.d(\wb_csr_data~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[8]~q ),
	.prn(vcc));
defparam \wb_csr_data[8] .is_wysiwyg = "true";
defparam \wb_csr_data[8] .power_up = "low";

cyclone10lp_lcell_comb \npc[8]~12 (
	.dataa(\pc_cntr[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[7]~11 ),
	.combout(\npc[8]~12_combout ),
	.cout(\npc[8]~13 ));
defparam \npc[8]~12 .lut_mask = 16'hA50A;
defparam \npc[8]~12 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~6 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[8]~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~6_combout ),
	.cout());
defparam \id_npc~6 .lut_mask = 16'h8080;
defparam \id_npc~6 .sum_lutc_input = "datac";

dffeas \id_npc[8] (
	.clk(clk_clk),
	.d(\id_npc~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[8]~q ),
	.prn(vcc));
defparam \id_npc[8] .is_wysiwyg = "true";
defparam \id_npc[8] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~6 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[8]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~6_combout ),
	.cout());
defparam \ex_npc~6 .lut_mask = 16'h8080;
defparam \ex_npc~6 .sum_lutc_input = "datac";

dffeas \ex_npc[8] (
	.clk(clk_clk),
	.d(\ex_npc~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[8]~q ),
	.prn(vcc));
defparam \ex_npc[8] .is_wysiwyg = "true";
defparam \ex_npc[8] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~4 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~4_combout ),
	.cout());
defparam \mem_npc~4 .lut_mask = 16'h8888;
defparam \mem_npc~4 .sum_lutc_input = "datac";

dffeas \mem_npc[8] (
	.clk(clk_clk),
	.d(\mem_npc~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[8]~q ),
	.prn(vcc));
defparam \mem_npc[8] .is_wysiwyg = "true";
defparam \mem_npc[8] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~4 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~4_combout ),
	.cout());
defparam \wb_npc~4 .lut_mask = 16'h8888;
defparam \wb_npc~4 .sum_lutc_input = "datac";

dffeas \wb_npc[8] (
	.clk(clk_clk),
	.d(\wb_npc~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[8]~q ),
	.prn(vcc));
defparam \wb_npc[8] .is_wysiwyg = "true";
defparam \wb_npc[8] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~6 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~6_combout ),
	.cout());
defparam \wb_alu_out~6 .lut_mask = 16'h8888;
defparam \wb_alu_out~6 .sum_lutc_input = "datac";

dffeas \wb_alu_out[8] (
	.clk(clk_clk),
	.d(\wb_alu_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[8]~q ),
	.prn(vcc));
defparam \wb_alu_out[8] .is_wysiwyg = "true";
defparam \wb_alu_out[8] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[8]~15 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[8]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[8]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[8]~15_combout ),
	.cout());
defparam \_T_3543__T_3854_data[8]~15 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[8]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[22]~89 (
	.dataa(mem_alu_out_0),
	.datab(mem_alu_out_1),
	.datac(Equal68),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_dmem_read_data[22]~89_combout ),
	.cout());
defparam \wb_dmem_read_data[22]~89 .lut_mask = 16'hB0B0;
defparam \wb_dmem_read_data[22]~89 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[22]~90 (
	.dataa(mem_alu_out_0),
	.datab(mem_alu_out_1),
	.datac(Equal68),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_dmem_read_data[22]~90_combout ),
	.cout());
defparam \wb_dmem_read_data[22]~90 .lut_mask = 16'hE0E0;
defparam \wb_dmem_read_data[22]~90 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~22 (
	.dataa(av_readdata_pre_24),
	.datab(av_readdata_pre_8),
	.datac(gnd),
	.datad(mem_alu_out_1),
	.cin(gnd),
	.combout(\wb_dmem_read_data~22_combout ),
	.cout());
defparam \wb_dmem_read_data~22 .lut_mask = 16'hAACC;
defparam \wb_dmem_read_data~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~43 (
	.dataa(\wb_dmem_read_data[22]~89_combout ),
	.datab(av_readdata_pre_23),
	.datac(\wb_dmem_read_data[22]~90_combout ),
	.datad(\wb_dmem_read_data~22_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~43_combout ),
	.cout());
defparam \wb_dmem_read_data~43 .lut_mask = 16'hE5E0;
defparam \wb_dmem_read_data~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~44 (
	.dataa(av_readdata_pre_7),
	.datab(\wb_dmem_read_data[22]~89_combout ),
	.datac(\wb_dmem_read_data~43_combout ),
	.datad(\wb_dmem_read_data~28_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~44_combout ),
	.cout());
defparam \wb_dmem_read_data~44 .lut_mask = 16'hF838;
defparam \wb_dmem_read_data~44 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[14]~45 (
	.dataa(\mem_ctrl_mask_type[0]~q ),
	.datab(\mem_ctrl_mask_type[1]~q ),
	.datac(gnd),
	.datad(mem_ctrl_mem_wr01),
	.cin(gnd),
	.combout(\wb_dmem_read_data[14]~45_combout ),
	.cout());
defparam \wb_dmem_read_data[14]~45 .lut_mask = 16'h99FF;
defparam \wb_dmem_read_data[14]~45 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[14]~46 (
	.dataa(mem_ctrl_mem_wr01),
	.datab(mem_alu_out_0),
	.datac(\mem_ctrl_mask_type[0]~q ),
	.datad(\mem_ctrl_mask_type[1]~q ),
	.cin(gnd),
	.combout(\wb_dmem_read_data[14]~46_combout ),
	.cout());
defparam \wb_dmem_read_data[14]~46 .lut_mask = 16'h08A0;
defparam \wb_dmem_read_data[14]~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[14]~47 (
	.dataa(\wb_dmem_read_data[14]~46_combout ),
	.datab(\wb_dmem_read_data[22]~90_combout ),
	.datac(\wb_dmem_read_data[22]~89_combout ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\wb_dmem_read_data[14]~47_combout ),
	.cout());
defparam \wb_dmem_read_data[14]~47 .lut_mask = 16'h02FF;
defparam \wb_dmem_read_data[14]~47 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~48 (
	.dataa(av_readdata_pre_8),
	.datab(\wb_dmem_read_data~44_combout ),
	.datac(\wb_dmem_read_data[14]~45_combout ),
	.datad(\wb_dmem_read_data[14]~47_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~48_combout ),
	.cout());
defparam \wb_dmem_read_data~48 .lut_mask = 16'h00AC;
defparam \wb_dmem_read_data~48 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[8] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[8]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[8] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[8] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[8]~16 (
	.dataa(\wb_csr_data[8]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[8]~15_combout ),
	.datad(\wb_dmem_read_data[8]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[8]~16_combout ),
	.cout());
defparam \_T_3543__T_3854_data[8]~16 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[8]~16 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a24 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[8]~16_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a24_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_a_first_bit_number = 24;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_b_first_bit_number = 24;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a24 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~9 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a24~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~9_combout ),
	.cout());
defparam \ex_rs_1~9 .lut_mask = 16'h8888;
defparam \ex_rs_1~9 .sum_lutc_input = "datac";

dffeas \ex_rs_1[8] (
	.clk(clk_clk),
	.d(\ex_rs_1~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[8]~q ),
	.prn(vcc));
defparam \ex_rs_1[8] .is_wysiwyg = "true";
defparam \ex_rs_1[8] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[8]~34 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_8),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[8]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[8]~34_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[8]~34 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[8]~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[8]~35 (
	.dataa(\ex_rs_1[8]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[8]~34_combout ),
	.datad(\wb_csr_data[8]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[8]~35_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[8]~35 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[8]~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[8]~36 (
	.dataa(\mem_alu_out[8]~q ),
	.datab(\ex_reg_rs2_bypass[8]~35_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[8]~36_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[8]~36 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[8]~36 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[8]~46 (
	.dataa(\_T_3681~3_combout ),
	.datab(\mem_csr_data[8]~q ),
	.datac(\ex_reg_rs2_bypass[8]~36_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\alu_io_op2[8]~46_combout ),
	.cout());
defparam \alu_io_op2[8]~46 .lut_mask = 16'hF8F8;
defparam \alu_io_op2[8]~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[8]~47 (
	.dataa(\alu_io_op2[5]~43_combout ),
	.datab(\ex_csr_addr[8]~q ),
	.datac(\ex_ctrl_alu_op2.10~q ),
	.datad(\alu_io_op2[8]~46_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[8]~47_combout ),
	.cout());
defparam \alu_io_op2[8]~47 .lut_mask = 16'hA808;
defparam \alu_io_op2[8]~47 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[8]~34 (
	.dataa(\ex_reg_rs1_bypass[0]~20_combout ),
	.datab(\mem_alu_out[8]~q ),
	.datac(\_T_3634~2_combout ),
	.datad(\mem_csr_data[8]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[8]~34_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[8]~34 .lut_mask = 16'hF888;
defparam \ex_reg_rs1_bypass[8]~34 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a24 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[8]~16_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a24_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_a_first_bit_number = 24;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_b_first_bit_number = 24;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a24 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~8 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a24~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~8_combout ),
	.cout());
defparam \ex_rs_0~8 .lut_mask = 16'h0080;
defparam \ex_rs_0~8 .sum_lutc_input = "datac";

dffeas \ex_rs_0[8] (
	.clk(clk_clk),
	.d(\ex_rs_0~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[8]~q ),
	.prn(vcc));
defparam \ex_rs_0[8] .is_wysiwyg = "true";
defparam \ex_rs_0[8] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[8]~35 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(av_readdata_pre_8),
	.datac(\wb_alu_out[8]~q ),
	.datad(\ex_reg_rs1_bypass[2]~138_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[8]~35_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[8]~35 .lut_mask = 16'hAAD8;
defparam \ex_reg_rs1_bypass[8]~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[8]~36 (
	.dataa(\ex_rs_0[8]~q ),
	.datab(\wb_csr_data[8]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\ex_reg_rs1_bypass[8]~35_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[8]~36_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[8]~36 .lut_mask = 16'hCFA0;
defparam \ex_reg_rs1_bypass[8]~36 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[8]~37 (
	.dataa(\ex_reg_rs1_bypass[0]~4_combout ),
	.datab(\ex_reg_rs1_bypass[8]~34_combout ),
	.datac(\ex_reg_rs1_bypass[8]~36_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[8]~37_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[8]~37 .lut_mask = 16'hECEC;
defparam \ex_reg_rs1_bypass[8]~37 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[8]~94 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[8]~q ),
	.datad(\ex_reg_rs1_bypass[8]~37_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[8]~94_combout ),
	.cout());
defparam \alu_io_op1[8]~94 .lut_mask = 16'h6240;
defparam \alu_io_op1[8]~94 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~155 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\alu_io_op2[8]~47_combout ),
	.datad(\alu_io_op1[8]~94_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~155_combout ),
	.cout());
defparam \mem_alu_out~155 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~155 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~156 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~155_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~173_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~156_combout ),
	.cout());
defparam \mem_alu_out~156 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~156 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~37 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[8]~94_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~156_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~37_combout ),
	.cout());
defparam \mem_alu_out~37 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~37 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~38 (
	.dataa(\alu_io_op2[8]~47_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~37_combout ),
	.datad(\alu|ShiftRight0~175_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~38_combout ),
	.cout());
defparam \mem_alu_out~38 .lut_mask = 16'hF838;
defparam \mem_alu_out~38 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~39 (
	.dataa(\mem_alu_out~38_combout ),
	.datab(\alu|_T_3[8]~16_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~39_combout ),
	.cout());
defparam \mem_alu_out~39 .lut_mask = 16'h00AC;
defparam \mem_alu_out~39 .sum_lutc_input = "datac";

dffeas \mem_alu_out[8] (
	.clk(clk_clk),
	.d(\mem_alu_out~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[8]~q ),
	.prn(vcc));
defparam \mem_alu_out[8] .is_wysiwyg = "true";
defparam \mem_alu_out[8] .power_up = "low";

cyclone10lp_lcell_comb \pc_cntr~28 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(\mem_alu_out[8]~q ),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[8]~12_combout ),
	.cin(gnd),
	.combout(\pc_cntr~28_combout ),
	.cout());
defparam \pc_cntr~28 .lut_mask = 16'hDAD0;
defparam \pc_cntr~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~29 (
	.dataa(\_T_3862[8]~16_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~28_combout ),
	.datad(\csr|mepc[8]~q ),
	.cin(gnd),
	.combout(\pc_cntr~29_combout ),
	.cout());
defparam \pc_cntr~29 .lut_mask = 16'hF2C2;
defparam \pc_cntr~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~30 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~29_combout ),
	.datac(\csr|mtvec[8]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~30_combout ),
	.cout());
defparam \pc_cntr~30 .lut_mask = 16'h88A0;
defparam \pc_cntr~30 .sum_lutc_input = "datac";

dffeas \pc_cntr[8] (
	.clk(clk_clk),
	.d(\pc_cntr~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[8]~q ),
	.prn(vcc));
defparam \pc_cntr[8] .is_wysiwyg = "true";
defparam \pc_cntr[8] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~7 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[8]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~7_combout ),
	.cout());
defparam \id_pc~7 .lut_mask = 16'h8080;
defparam \id_pc~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~7 (
	.dataa(id_pc_9),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~7_combout ),
	.cout());
defparam \ex_pc~7 .lut_mask = 16'h8080;
defparam \ex_pc~7 .sum_lutc_input = "datac";

dffeas \ex_pc[9] (
	.clk(clk_clk),
	.d(\ex_pc~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[9]~q ),
	.prn(vcc));
defparam \ex_pc[9] .is_wysiwyg = "true";
defparam \ex_pc[9] .power_up = "low";

cyclone10lp_lcell_comb \mem_csr_data~14 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[9]~66_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~14_combout ),
	.cout());
defparam \mem_csr_data~14 .lut_mask = 16'h8888;
defparam \mem_csr_data~14 .sum_lutc_input = "datac";

dffeas \mem_csr_data[9] (
	.clk(clk_clk),
	.d(\mem_csr_data~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[9]~q ),
	.prn(vcc));
defparam \mem_csr_data[9] .is_wysiwyg = "true";
defparam \mem_csr_data[9] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[9]~38 (
	.dataa(\ex_reg_rs1_bypass[0]~20_combout ),
	.datab(\mem_alu_out[9]~q ),
	.datac(\_T_3634~2_combout ),
	.datad(\mem_csr_data[9]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[9]~38_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[9]~38 .lut_mask = 16'hF888;
defparam \ex_reg_rs1_bypass[9]~38 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_csr_data~7 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~7_combout ),
	.cout());
defparam \wb_csr_data~7 .lut_mask = 16'h8888;
defparam \wb_csr_data~7 .sum_lutc_input = "datac";

dffeas \wb_csr_data[9] (
	.clk(clk_clk),
	.d(\wb_csr_data~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[9]~q ),
	.prn(vcc));
defparam \wb_csr_data[9] .is_wysiwyg = "true";
defparam \wb_csr_data[9] .power_up = "low";

cyclone10lp_lcell_comb \npc[9]~14 (
	.dataa(\pc_cntr[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[8]~13 ),
	.combout(\npc[9]~14_combout ),
	.cout(\npc[9]~15 ));
defparam \npc[9]~14 .lut_mask = 16'h5A5F;
defparam \npc[9]~14 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~7 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[9]~14_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~7_combout ),
	.cout());
defparam \id_npc~7 .lut_mask = 16'h8080;
defparam \id_npc~7 .sum_lutc_input = "datac";

dffeas \id_npc[9] (
	.clk(clk_clk),
	.d(\id_npc~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[9]~q ),
	.prn(vcc));
defparam \id_npc[9] .is_wysiwyg = "true";
defparam \id_npc[9] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~7 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~7_combout ),
	.cout());
defparam \ex_npc~7 .lut_mask = 16'h8080;
defparam \ex_npc~7 .sum_lutc_input = "datac";

dffeas \ex_npc[9] (
	.clk(clk_clk),
	.d(\ex_npc~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[9]~q ),
	.prn(vcc));
defparam \ex_npc[9] .is_wysiwyg = "true";
defparam \ex_npc[9] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~5 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~5_combout ),
	.cout());
defparam \mem_npc~5 .lut_mask = 16'h8888;
defparam \mem_npc~5 .sum_lutc_input = "datac";

dffeas \mem_npc[9] (
	.clk(clk_clk),
	.d(\mem_npc~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[9]~q ),
	.prn(vcc));
defparam \mem_npc[9] .is_wysiwyg = "true";
defparam \mem_npc[9] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~5 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~5_combout ),
	.cout());
defparam \wb_npc~5 .lut_mask = 16'h8888;
defparam \wb_npc~5 .sum_lutc_input = "datac";

dffeas \wb_npc[9] (
	.clk(clk_clk),
	.d(\wb_npc~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[9]~q ),
	.prn(vcc));
defparam \wb_npc[9] .is_wysiwyg = "true";
defparam \wb_npc[9] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~7 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~7_combout ),
	.cout());
defparam \wb_alu_out~7 .lut_mask = 16'h8888;
defparam \wb_alu_out~7 .sum_lutc_input = "datac";

dffeas \wb_alu_out[9] (
	.clk(clk_clk),
	.d(\wb_alu_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[9]~q ),
	.prn(vcc));
defparam \wb_alu_out[9] .is_wysiwyg = "true";
defparam \wb_alu_out[9] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[9]~17 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[9]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[9]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[9]~17_combout ),
	.cout());
defparam \_T_3543__T_3854_data[9]~17 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[9]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~16 (
	.dataa(av_readdata_pre_25),
	.datab(av_readdata_pre_9),
	.datac(gnd),
	.datad(mem_alu_out_1),
	.cin(gnd),
	.combout(\wb_dmem_read_data~16_combout ),
	.cout());
defparam \wb_dmem_read_data~16 .lut_mask = 16'hAACC;
defparam \wb_dmem_read_data~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~49 (
	.dataa(\wb_dmem_read_data[22]~90_combout ),
	.datab(av_readdata_pre_7),
	.datac(\wb_dmem_read_data[22]~89_combout ),
	.datad(\wb_dmem_read_data~16_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~49_combout ),
	.cout());
defparam \wb_dmem_read_data~49 .lut_mask = 16'hE5E0;
defparam \wb_dmem_read_data~49 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~50 (
	.dataa(av_readdata_pre_23),
	.datab(\wb_dmem_read_data[22]~90_combout ),
	.datac(\wb_dmem_read_data~49_combout ),
	.datad(\wb_dmem_read_data~28_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~50_combout ),
	.cout());
defparam \wb_dmem_read_data~50 .lut_mask = 16'hF838;
defparam \wb_dmem_read_data~50 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~51 (
	.dataa(av_readdata_pre_9),
	.datab(\wb_dmem_read_data~50_combout ),
	.datac(\wb_dmem_read_data[14]~45_combout ),
	.datad(\wb_dmem_read_data[14]~47_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~51_combout ),
	.cout());
defparam \wb_dmem_read_data~51 .lut_mask = 16'h00AC;
defparam \wb_dmem_read_data~51 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[9] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[9]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[9] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[9] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[9]~18 (
	.dataa(\wb_npc[9]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[9]~17_combout ),
	.datad(\wb_dmem_read_data[9]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[9]~18_combout ),
	.cout());
defparam \_T_3543__T_3854_data[9]~18 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[9]~18 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a23 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[9]~18_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a23_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_a_first_bit_number = 23;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_b_first_bit_number = 23;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a23 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~9 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a23~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~9_combout ),
	.cout());
defparam \ex_rs_0~9 .lut_mask = 16'h0080;
defparam \ex_rs_0~9 .sum_lutc_input = "datac";

dffeas \ex_rs_0[9] (
	.clk(clk_clk),
	.d(\ex_rs_0~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[9]~q ),
	.prn(vcc));
defparam \ex_rs_0[9] .is_wysiwyg = "true";
defparam \ex_rs_0[9] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[9]~39 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(\ex_rs_0[9]~q ),
	.datac(\wb_alu_out[9]~q ),
	.datad(\ex_reg_rs1_bypass[2]~7_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[9]~39_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[9]~39 .lut_mask = 16'hAAD8;
defparam \ex_reg_rs1_bypass[9]~39 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[9]~40 (
	.dataa(av_readdata_pre_9),
	.datab(\wb_csr_data[9]~q ),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\ex_reg_rs1_bypass[9]~39_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[9]~40_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[9]~40 .lut_mask = 16'hCFA0;
defparam \ex_reg_rs1_bypass[9]~40 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[9]~41 (
	.dataa(\ex_reg_rs1_bypass[0]~4_combout ),
	.datab(\ex_reg_rs1_bypass[9]~38_combout ),
	.datac(\ex_reg_rs1_bypass[9]~40_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[9]~41_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[9]~41 .lut_mask = 16'hECEC;
defparam \ex_reg_rs1_bypass[9]~41 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[9]~95 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[9]~q ),
	.datad(\ex_reg_rs1_bypass[9]~41_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[9]~95_combout ),
	.cout());
defparam \alu_io_op1[9]~95 .lut_mask = 16'h6240;
defparam \alu_io_op1[9]~95 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_csr_addr~6 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[29]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_csr_addr~6_combout ),
	.cout());
defparam \ex_csr_addr~6 .lut_mask = 16'h8080;
defparam \ex_csr_addr~6 .sum_lutc_input = "datac";

dffeas \ex_csr_addr[9] (
	.clk(clk_clk),
	.d(\ex_csr_addr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_addr[9]~q ),
	.prn(vcc));
defparam \ex_csr_addr[9] .is_wysiwyg = "true";
defparam \ex_csr_addr[9] .power_up = "low";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a23 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[9]~18_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a23_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_a_first_bit_number = 23;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_b_first_bit_number = 23;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a23 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~8 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a23~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~8_combout ),
	.cout());
defparam \ex_rs_1~8 .lut_mask = 16'h8888;
defparam \ex_rs_1~8 .sum_lutc_input = "datac";

dffeas \ex_rs_1[9] (
	.clk(clk_clk),
	.d(\ex_rs_1~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[9]~q ),
	.prn(vcc));
defparam \ex_rs_1[9] .is_wysiwyg = "true";
defparam \ex_rs_1[9] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[9]~31 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(\ex_rs_1[9]~q ),
	.datac(\wb_alu_out[9]~q ),
	.datad(\ex_reg_rs2_bypass[7]~5_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[9]~31_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[9]~31 .lut_mask = 16'hAAD8;
defparam \ex_reg_rs2_bypass[9]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[9]~32 (
	.dataa(av_readdata_pre_9),
	.datab(\wb_csr_data[9]~q ),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\ex_reg_rs2_bypass[9]~31_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[9]~32_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[9]~32 .lut_mask = 16'hCFA0;
defparam \ex_reg_rs2_bypass[9]~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[9]~33 (
	.dataa(\mem_alu_out[9]~q ),
	.datab(\_T_3686~0_combout ),
	.datac(\_T_3681~3_combout ),
	.datad(\ex_reg_rs2_bypass[9]~32_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[9]~33_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[9]~33 .lut_mask = 16'h0B08;
defparam \ex_reg_rs2_bypass[9]~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[9]~44 (
	.dataa(\_T_3681~3_combout ),
	.datab(\mem_csr_data[9]~q ),
	.datac(\ex_reg_rs2_bypass[9]~33_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\alu_io_op2[9]~44_combout ),
	.cout());
defparam \alu_io_op2[9]~44 .lut_mask = 16'hF8F8;
defparam \alu_io_op2[9]~44 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[9]~45 (
	.dataa(\alu_io_op2[5]~43_combout ),
	.datab(\ex_csr_addr[9]~q ),
	.datac(\ex_ctrl_alu_op2.10~q ),
	.datad(\alu_io_op2[9]~44_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[9]~45_combout ),
	.cout());
defparam \alu_io_op2[9]~45 .lut_mask = 16'hA808;
defparam \alu_io_op2[9]~45 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~153 (
	.dataa(\mem_alu_out[26]~2_combout ),
	.datab(\alu|LessThan0~0_combout ),
	.datac(\alu_io_op2[9]~45_combout ),
	.datad(\alu_io_op1[9]~95_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~153_combout ),
	.cout());
defparam \mem_alu_out~153 .lut_mask = 16'h7DD4;
defparam \mem_alu_out~153 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~154 (
	.dataa(\mem_alu_out[26]~2_combout ),
	.datab(\mem_alu_out~153_combout ),
	.datac(\alu|LessThan0~0_combout ),
	.datad(\alu|ShiftRight0~180_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~154_combout ),
	.cout());
defparam \mem_alu_out~154 .lut_mask = 16'hCC8C;
defparam \mem_alu_out~154 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~40 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[9]~45_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~154_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~40_combout ),
	.cout());
defparam \mem_alu_out~40 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~40 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~41 (
	.dataa(\alu_io_op1[9]~95_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~40_combout ),
	.datad(\alu|ShiftRight0~183_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~41_combout ),
	.cout());
defparam \mem_alu_out~41 .lut_mask = 16'hF838;
defparam \mem_alu_out~41 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~42 (
	.dataa(\mem_alu_out~41_combout ),
	.datab(\alu|_T_3[9]~18_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~42_combout ),
	.cout());
defparam \mem_alu_out~42 .lut_mask = 16'h00AC;
defparam \mem_alu_out~42 .sum_lutc_input = "datac";

dffeas \mem_alu_out[9] (
	.clk(clk_clk),
	.d(\mem_alu_out~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[9]~q ),
	.prn(vcc));
defparam \mem_alu_out[9] .is_wysiwyg = "true";
defparam \mem_alu_out[9] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~7 (
	.dataa(\ex_pc[9]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~7_combout ),
	.cout());
defparam \mem_pc~7 .lut_mask = 16'h8888;
defparam \mem_pc~7 .sum_lutc_input = "datac";

dffeas \mem_pc[9] (
	.clk(clk_clk),
	.d(\mem_pc~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[9]~q ),
	.prn(vcc));
defparam \mem_pc[9] .is_wysiwyg = "true";
defparam \mem_pc[9] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~24 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_csr_addr[9]~q ),
	.datac(\ex_ctrl_imm_type.101~q ),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\mem_imm~24_combout ),
	.cout());
defparam \mem_imm~24 .lut_mask = 16'h0008;
defparam \mem_imm~24 .sum_lutc_input = "datac";

dffeas \mem_imm[9] (
	.clk(clk_clk),
	.d(\mem_imm~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[9]~q ),
	.prn(vcc));
defparam \mem_imm[9] .is_wysiwyg = "true";
defparam \mem_imm[9] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[9]~18 (
	.dataa(\mem_pc[9]~q ),
	.datab(\mem_imm[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[8]~17 ),
	.combout(\_T_3862[9]~18_combout ),
	.cout(\_T_3862[9]~19 ));
defparam \_T_3862[9]~18 .lut_mask = 16'h9617;
defparam \_T_3862[9]~18 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~31 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[9]~18_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[9]~14_combout ),
	.cin(gnd),
	.combout(\pc_cntr~31_combout ),
	.cout());
defparam \pc_cntr~31 .lut_mask = 16'h5E0E;
defparam \pc_cntr~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~32 (
	.dataa(\mem_alu_out[9]~q ),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~31_combout ),
	.datad(\csr|mepc[9]~q ),
	.cin(gnd),
	.combout(\pc_cntr~32_combout ),
	.cout());
defparam \pc_cntr~32 .lut_mask = 16'hF838;
defparam \pc_cntr~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~33 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~32_combout ),
	.datac(\csr|mtvec[9]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~33_combout ),
	.cout());
defparam \pc_cntr~33 .lut_mask = 16'h88A0;
defparam \pc_cntr~33 .sum_lutc_input = "datac";

dffeas \pc_cntr[9] (
	.clk(clk_clk),
	.d(\pc_cntr~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[9]~q ),
	.prn(vcc));
defparam \pc_cntr[9] .is_wysiwyg = "true";
defparam \pc_cntr[9] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~8 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~8_combout ),
	.cout());
defparam \id_pc~8 .lut_mask = 16'h8080;
defparam \id_pc~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~8 (
	.dataa(id_pc_10),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~8_combout ),
	.cout());
defparam \ex_pc~8 .lut_mask = 16'h8080;
defparam \ex_pc~8 .sum_lutc_input = "datac";

dffeas \ex_pc[10] (
	.clk(clk_clk),
	.d(\ex_pc~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[10]~q ),
	.prn(vcc));
defparam \ex_pc[10] .is_wysiwyg = "true";
defparam \ex_pc[10] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~8 (
	.dataa(\ex_pc[10]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~8_combout ),
	.cout());
defparam \mem_pc~8 .lut_mask = 16'h8888;
defparam \mem_pc~8 .sum_lutc_input = "datac";

dffeas \mem_pc[10] (
	.clk(clk_clk),
	.d(\mem_pc~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[10]~q ),
	.prn(vcc));
defparam \mem_pc[10] .is_wysiwyg = "true";
defparam \mem_pc[10] .power_up = "low";

cyclone10lp_lcell_comb \ex_csr_addr~8 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[30]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_csr_addr~8_combout ),
	.cout());
defparam \ex_csr_addr~8 .lut_mask = 16'h8080;
defparam \ex_csr_addr~8 .sum_lutc_input = "datac";

dffeas \ex_csr_addr[10] (
	.clk(clk_clk),
	.d(\ex_csr_addr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_addr[10]~q ),
	.prn(vcc));
defparam \ex_csr_addr[10] .is_wysiwyg = "true";
defparam \ex_csr_addr[10] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~25 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_csr_addr[10]~q ),
	.datac(\ex_ctrl_imm_type.101~q ),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\mem_imm~25_combout ),
	.cout());
defparam \mem_imm~25 .lut_mask = 16'h0008;
defparam \mem_imm~25 .sum_lutc_input = "datac";

dffeas \mem_imm[10] (
	.clk(clk_clk),
	.d(\mem_imm~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[10]~q ),
	.prn(vcc));
defparam \mem_imm[10] .is_wysiwyg = "true";
defparam \mem_imm[10] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[10]~20 (
	.dataa(\mem_pc[10]~q ),
	.datab(\mem_imm[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[9]~19 ),
	.combout(\_T_3862[10]~20_combout ),
	.cout(\_T_3862[10]~21 ));
defparam \_T_3862[10]~20 .lut_mask = 16'h698E;
defparam \_T_3862[10]~20 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \mem_csr_data~15 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[10]~72_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~15_combout ),
	.cout());
defparam \mem_csr_data~15 .lut_mask = 16'h8888;
defparam \mem_csr_data~15 .sum_lutc_input = "datac";

dffeas \mem_csr_data[10] (
	.clk(clk_clk),
	.d(\mem_csr_data~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[10]~q ),
	.prn(vcc));
defparam \mem_csr_data[10] .is_wysiwyg = "true";
defparam \mem_csr_data[10] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~8 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~8_combout ),
	.cout());
defparam \wb_csr_data~8 .lut_mask = 16'h8888;
defparam \wb_csr_data~8 .sum_lutc_input = "datac";

dffeas \wb_csr_data[10] (
	.clk(clk_clk),
	.d(\wb_csr_data~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[10]~q ),
	.prn(vcc));
defparam \wb_csr_data[10] .is_wysiwyg = "true";
defparam \wb_csr_data[10] .power_up = "low";

cyclone10lp_lcell_comb \npc[10]~16 (
	.dataa(\pc_cntr[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[9]~15 ),
	.combout(\npc[10]~16_combout ),
	.cout(\npc[10]~17 ));
defparam \npc[10]~16 .lut_mask = 16'hA50A;
defparam \npc[10]~16 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~8 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[10]~16_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~8_combout ),
	.cout());
defparam \id_npc~8 .lut_mask = 16'h8080;
defparam \id_npc~8 .sum_lutc_input = "datac";

dffeas \id_npc[10] (
	.clk(clk_clk),
	.d(\id_npc~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[10]~q ),
	.prn(vcc));
defparam \id_npc[10] .is_wysiwyg = "true";
defparam \id_npc[10] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~8 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[10]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~8_combout ),
	.cout());
defparam \ex_npc~8 .lut_mask = 16'h8080;
defparam \ex_npc~8 .sum_lutc_input = "datac";

dffeas \ex_npc[10] (
	.clk(clk_clk),
	.d(\ex_npc~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[10]~q ),
	.prn(vcc));
defparam \ex_npc[10] .is_wysiwyg = "true";
defparam \ex_npc[10] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~6 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~6_combout ),
	.cout());
defparam \mem_npc~6 .lut_mask = 16'h8888;
defparam \mem_npc~6 .sum_lutc_input = "datac";

dffeas \mem_npc[10] (
	.clk(clk_clk),
	.d(\mem_npc~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[10]~q ),
	.prn(vcc));
defparam \mem_npc[10] .is_wysiwyg = "true";
defparam \mem_npc[10] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~6 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~6_combout ),
	.cout());
defparam \wb_npc~6 .lut_mask = 16'h8888;
defparam \wb_npc~6 .sum_lutc_input = "datac";

dffeas \wb_npc[10] (
	.clk(clk_clk),
	.d(\wb_npc~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[10]~q ),
	.prn(vcc));
defparam \wb_npc[10] .is_wysiwyg = "true";
defparam \wb_npc[10] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~8 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~8_combout ),
	.cout());
defparam \wb_alu_out~8 .lut_mask = 16'h8888;
defparam \wb_alu_out~8 .sum_lutc_input = "datac";

dffeas \wb_alu_out[10] (
	.clk(clk_clk),
	.d(\wb_alu_out~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[10]~q ),
	.prn(vcc));
defparam \wb_alu_out[10] .is_wysiwyg = "true";
defparam \wb_alu_out[10] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[10]~19 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[10]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[10]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[10]~19_combout ),
	.cout());
defparam \_T_3543__T_3854_data[10]~19 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[10]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~52 (
	.dataa(av_readdata_pre_26),
	.datab(av_readdata_pre_10),
	.datac(gnd),
	.datad(mem_alu_out_1),
	.cin(gnd),
	.combout(\wb_dmem_read_data~52_combout ),
	.cout());
defparam \wb_dmem_read_data~52 .lut_mask = 16'hAACC;
defparam \wb_dmem_read_data~52 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~53 (
	.dataa(\wb_dmem_read_data[22]~89_combout ),
	.datab(av_readdata_pre_23),
	.datac(\wb_dmem_read_data[22]~90_combout ),
	.datad(\wb_dmem_read_data~52_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~53_combout ),
	.cout());
defparam \wb_dmem_read_data~53 .lut_mask = 16'hE5E0;
defparam \wb_dmem_read_data~53 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~54 (
	.dataa(av_readdata_pre_7),
	.datab(\wb_dmem_read_data[22]~89_combout ),
	.datac(\wb_dmem_read_data~53_combout ),
	.datad(\wb_dmem_read_data~28_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~54_combout ),
	.cout());
defparam \wb_dmem_read_data~54 .lut_mask = 16'hF838;
defparam \wb_dmem_read_data~54 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~55 (
	.dataa(av_readdata_pre_10),
	.datab(\wb_dmem_read_data~54_combout ),
	.datac(\wb_dmem_read_data[14]~45_combout ),
	.datad(\wb_dmem_read_data[14]~47_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~55_combout ),
	.cout());
defparam \wb_dmem_read_data~55 .lut_mask = 16'h00AC;
defparam \wb_dmem_read_data~55 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[10] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[10]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[10] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[10] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[10]~20 (
	.dataa(\wb_csr_data[10]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[10]~19_combout ),
	.datad(\wb_dmem_read_data[10]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[10]~20_combout ),
	.cout());
defparam \_T_3543__T_3854_data[10]~20 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[10]~20 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a22 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[10]~20_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a22_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_a_first_bit_number = 22;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_b_first_bit_number = 22;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a22 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~10 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a22~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~10_combout ),
	.cout());
defparam \ex_rs_1~10 .lut_mask = 16'h8888;
defparam \ex_rs_1~10 .sum_lutc_input = "datac";

dffeas \ex_rs_1[10] (
	.clk(clk_clk),
	.d(\ex_rs_1~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[10]~q ),
	.prn(vcc));
defparam \ex_rs_1[10] .is_wysiwyg = "true";
defparam \ex_rs_1[10] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[10]~37 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_10),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[10]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[10]~37_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[10]~37 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[10]~37 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[10]~38 (
	.dataa(\ex_rs_1[10]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[10]~37_combout ),
	.datad(\wb_csr_data[10]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[10]~38_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[10]~38 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[10]~38 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[10]~39 (
	.dataa(\mem_alu_out[10]~q ),
	.datab(\ex_reg_rs2_bypass[10]~38_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[10]~39_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[10]~39 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[10]~39 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[10]~48 (
	.dataa(\_T_3681~3_combout ),
	.datab(\mem_csr_data[10]~q ),
	.datac(\ex_reg_rs2_bypass[10]~39_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\alu_io_op2[10]~48_combout ),
	.cout());
defparam \alu_io_op2[10]~48 .lut_mask = 16'hF8F8;
defparam \alu_io_op2[10]~48 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[10]~49 (
	.dataa(\alu_io_op2[5]~43_combout ),
	.datab(\ex_csr_addr[10]~q ),
	.datac(\ex_ctrl_alu_op2.10~q ),
	.datad(\alu_io_op2[10]~48_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[10]~49_combout ),
	.cout());
defparam \alu_io_op2[10]~49 .lut_mask = 16'hA808;
defparam \alu_io_op2[10]~49 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a22 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[10]~20_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a22_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_a_first_bit_number = 22;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_b_first_bit_number = 22;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a22 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~10 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a22~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~10_combout ),
	.cout());
defparam \ex_rs_0~10 .lut_mask = 16'h0080;
defparam \ex_rs_0~10 .sum_lutc_input = "datac";

dffeas \ex_rs_0[10] (
	.clk(clk_clk),
	.d(\ex_rs_0~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[10]~q ),
	.prn(vcc));
defparam \ex_rs_0[10] .is_wysiwyg = "true";
defparam \ex_rs_0[10] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[10]~42 (
	.dataa(\ex_rs_0[10]~q ),
	.datab(\wb_csr_data[10]~q ),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[10]~42_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[10]~42 .lut_mask = 16'hCACA;
defparam \ex_reg_rs1_bypass[10]~42 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[10]~43 (
	.dataa(av_readdata_pre_10),
	.datab(\ex_reg_rs1_bypass[2]~7_combout ),
	.datac(\wb_alu_out[10]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[10]~43_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[10]~43 .lut_mask = 16'hB8B8;
defparam \ex_reg_rs1_bypass[10]~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[10]~44 (
	.dataa(\ex_reg_rs1_bypass[0]~4_combout ),
	.datab(\ex_reg_rs1_bypass[2]~138_combout ),
	.datac(\ex_reg_rs1_bypass[10]~42_combout ),
	.datad(\ex_reg_rs1_bypass[10]~43_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[10]~44_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[10]~44 .lut_mask = 16'hA280;
defparam \ex_reg_rs1_bypass[10]~44 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[10]~139 (
	.dataa(\Equal59~0_combout ),
	.datab(\ex_inst[19]~q ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\mem_csr_data[10]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[10]~139_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[10]~139 .lut_mask = 16'hD000;
defparam \ex_reg_rs1_bypass[10]~139 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[10]~45 (
	.dataa(\ex_reg_rs1_bypass[0]~20_combout ),
	.datab(\mem_alu_out[10]~q ),
	.datac(\ex_reg_rs1_bypass[10]~44_combout ),
	.datad(\ex_reg_rs1_bypass[10]~139_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[10]~45_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[10]~45 .lut_mask = 16'hFFF8;
defparam \ex_reg_rs1_bypass[10]~45 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[10]~96 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[10]~q ),
	.datad(\ex_reg_rs1_bypass[10]~45_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[10]~96_combout ),
	.cout());
defparam \alu_io_op1[10]~96 .lut_mask = 16'h6240;
defparam \alu_io_op1[10]~96 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~151 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\alu_io_op2[10]~49_combout ),
	.datad(\alu_io_op1[10]~96_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~151_combout ),
	.cout());
defparam \mem_alu_out~151 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~151 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~152 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~151_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~188_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~152_combout ),
	.cout());
defparam \mem_alu_out~152 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~152 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~43 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[10]~96_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~152_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~43_combout ),
	.cout());
defparam \mem_alu_out~43 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~44 (
	.dataa(\alu_io_op2[10]~49_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~43_combout ),
	.datad(\alu|ShiftRight0~190_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~44_combout ),
	.cout());
defparam \mem_alu_out~44 .lut_mask = 16'hF838;
defparam \mem_alu_out~44 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~45 (
	.dataa(\mem_alu_out~44_combout ),
	.datab(\alu|_T_3[10]~20_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~45_combout ),
	.cout());
defparam \mem_alu_out~45 .lut_mask = 16'h00AC;
defparam \mem_alu_out~45 .sum_lutc_input = "datac";

dffeas \mem_alu_out[10] (
	.clk(clk_clk),
	.d(\mem_alu_out~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[10]~q ),
	.prn(vcc));
defparam \mem_alu_out[10] .is_wysiwyg = "true";
defparam \mem_alu_out[10] .power_up = "low";

cyclone10lp_lcell_comb \pc_cntr~34 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(\mem_alu_out[10]~q ),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[10]~16_combout ),
	.cin(gnd),
	.combout(\pc_cntr~34_combout ),
	.cout());
defparam \pc_cntr~34 .lut_mask = 16'hDAD0;
defparam \pc_cntr~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~35 (
	.dataa(\_T_3862[10]~20_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~34_combout ),
	.datad(\csr|mepc[10]~q ),
	.cin(gnd),
	.combout(\pc_cntr~35_combout ),
	.cout());
defparam \pc_cntr~35 .lut_mask = 16'hF2C2;
defparam \pc_cntr~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~36 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~35_combout ),
	.datac(\csr|mtvec[10]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~36_combout ),
	.cout());
defparam \pc_cntr~36 .lut_mask = 16'h88A0;
defparam \pc_cntr~36 .sum_lutc_input = "datac";

dffeas \pc_cntr[10] (
	.clk(clk_clk),
	.d(\pc_cntr~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[10]~q ),
	.prn(vcc));
defparam \pc_cntr[10] .is_wysiwyg = "true";
defparam \pc_cntr[10] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~9 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[10]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~9_combout ),
	.cout());
defparam \id_pc~9 .lut_mask = 16'h8080;
defparam \id_pc~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~9 (
	.dataa(id_pc_11),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~9_combout ),
	.cout());
defparam \ex_pc~9 .lut_mask = 16'h8080;
defparam \ex_pc~9 .sum_lutc_input = "datac";

dffeas \ex_pc[11] (
	.clk(clk_clk),
	.d(\ex_pc~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[11]~q ),
	.prn(vcc));
defparam \ex_pc[11] .is_wysiwyg = "true";
defparam \ex_pc[11] .power_up = "low";

cyclone10lp_lcell_comb \mem_csr_data~16 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[11]~79_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~16_combout ),
	.cout());
defparam \mem_csr_data~16 .lut_mask = 16'h8888;
defparam \mem_csr_data~16 .sum_lutc_input = "datac";

dffeas \mem_csr_data[11] (
	.clk(clk_clk),
	.d(\mem_csr_data~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[11]~q ),
	.prn(vcc));
defparam \mem_csr_data[11] .is_wysiwyg = "true";
defparam \mem_csr_data[11] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[11]~46 (
	.dataa(\ex_reg_rs1_bypass[0]~20_combout ),
	.datab(\mem_alu_out[11]~q ),
	.datac(\_T_3634~2_combout ),
	.datad(\mem_csr_data[11]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[11]~46_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[11]~46 .lut_mask = 16'hF888;
defparam \ex_reg_rs1_bypass[11]~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_csr_data~9 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~9_combout ),
	.cout());
defparam \wb_csr_data~9 .lut_mask = 16'h8888;
defparam \wb_csr_data~9 .sum_lutc_input = "datac";

dffeas \wb_csr_data[11] (
	.clk(clk_clk),
	.d(\wb_csr_data~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[11]~q ),
	.prn(vcc));
defparam \wb_csr_data[11] .is_wysiwyg = "true";
defparam \wb_csr_data[11] .power_up = "low";

cyclone10lp_lcell_comb \npc[11]~18 (
	.dataa(\pc_cntr[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[10]~17 ),
	.combout(\npc[11]~18_combout ),
	.cout(\npc[11]~19 ));
defparam \npc[11]~18 .lut_mask = 16'h5A5F;
defparam \npc[11]~18 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~9 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[11]~18_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~9_combout ),
	.cout());
defparam \id_npc~9 .lut_mask = 16'h8080;
defparam \id_npc~9 .sum_lutc_input = "datac";

dffeas \id_npc[11] (
	.clk(clk_clk),
	.d(\id_npc~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[11]~q ),
	.prn(vcc));
defparam \id_npc[11] .is_wysiwyg = "true";
defparam \id_npc[11] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~9 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[11]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~9_combout ),
	.cout());
defparam \ex_npc~9 .lut_mask = 16'h8080;
defparam \ex_npc~9 .sum_lutc_input = "datac";

dffeas \ex_npc[11] (
	.clk(clk_clk),
	.d(\ex_npc~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[11]~q ),
	.prn(vcc));
defparam \ex_npc[11] .is_wysiwyg = "true";
defparam \ex_npc[11] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~7 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~7_combout ),
	.cout());
defparam \mem_npc~7 .lut_mask = 16'h8888;
defparam \mem_npc~7 .sum_lutc_input = "datac";

dffeas \mem_npc[11] (
	.clk(clk_clk),
	.d(\mem_npc~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[11]~q ),
	.prn(vcc));
defparam \mem_npc[11] .is_wysiwyg = "true";
defparam \mem_npc[11] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~7 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~7_combout ),
	.cout());
defparam \wb_npc~7 .lut_mask = 16'h8888;
defparam \wb_npc~7 .sum_lutc_input = "datac";

dffeas \wb_npc[11] (
	.clk(clk_clk),
	.d(\wb_npc~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[11]~q ),
	.prn(vcc));
defparam \wb_npc[11] .is_wysiwyg = "true";
defparam \wb_npc[11] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~9 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~9_combout ),
	.cout());
defparam \wb_alu_out~9 .lut_mask = 16'h8888;
defparam \wb_alu_out~9 .sum_lutc_input = "datac";

dffeas \wb_alu_out[11] (
	.clk(clk_clk),
	.d(\wb_alu_out~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[11]~q ),
	.prn(vcc));
defparam \wb_alu_out[11] .is_wysiwyg = "true";
defparam \wb_alu_out[11] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[11]~21 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[11]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[11]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[11]~21_combout ),
	.cout());
defparam \_T_3543__T_3854_data[11]~21 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[11]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~56 (
	.dataa(av_readdata_pre_27),
	.datab(av_readdata_pre_11),
	.datac(gnd),
	.datad(mem_alu_out_1),
	.cin(gnd),
	.combout(\wb_dmem_read_data~56_combout ),
	.cout());
defparam \wb_dmem_read_data~56 .lut_mask = 16'hAACC;
defparam \wb_dmem_read_data~56 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~57 (
	.dataa(\wb_dmem_read_data[22]~90_combout ),
	.datab(av_readdata_pre_7),
	.datac(\wb_dmem_read_data[22]~89_combout ),
	.datad(\wb_dmem_read_data~56_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~57_combout ),
	.cout());
defparam \wb_dmem_read_data~57 .lut_mask = 16'hE5E0;
defparam \wb_dmem_read_data~57 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~58 (
	.dataa(av_readdata_pre_23),
	.datab(\wb_dmem_read_data[22]~90_combout ),
	.datac(\wb_dmem_read_data~57_combout ),
	.datad(\wb_dmem_read_data~28_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~58_combout ),
	.cout());
defparam \wb_dmem_read_data~58 .lut_mask = 16'hF838;
defparam \wb_dmem_read_data~58 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~59 (
	.dataa(av_readdata_pre_11),
	.datab(\wb_dmem_read_data~58_combout ),
	.datac(\wb_dmem_read_data[14]~45_combout ),
	.datad(\wb_dmem_read_data[14]~47_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~59_combout ),
	.cout());
defparam \wb_dmem_read_data~59 .lut_mask = 16'h00AC;
defparam \wb_dmem_read_data~59 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[11] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[11]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[11] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[11] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[11]~22 (
	.dataa(\wb_npc[11]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[11]~21_combout ),
	.datad(\wb_dmem_read_data[11]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[11]~22_combout ),
	.cout());
defparam \_T_3543__T_3854_data[11]~22 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[11]~22 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a21 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[11]~22_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a21_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_a_first_bit_number = 21;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_b_first_bit_number = 21;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a21 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~11 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a21~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~11_combout ),
	.cout());
defparam \ex_rs_0~11 .lut_mask = 16'h0080;
defparam \ex_rs_0~11 .sum_lutc_input = "datac";

dffeas \ex_rs_0[11] (
	.clk(clk_clk),
	.d(\ex_rs_0~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[11]~q ),
	.prn(vcc));
defparam \ex_rs_0[11] .is_wysiwyg = "true";
defparam \ex_rs_0[11] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[11]~47 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(\ex_rs_0[11]~q ),
	.datac(\wb_alu_out[11]~q ),
	.datad(\ex_reg_rs1_bypass[2]~7_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[11]~47_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[11]~47 .lut_mask = 16'hAAD8;
defparam \ex_reg_rs1_bypass[11]~47 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[11]~48 (
	.dataa(av_readdata_pre_11),
	.datab(\wb_csr_data[11]~q ),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\ex_reg_rs1_bypass[11]~47_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[11]~48_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[11]~48 .lut_mask = 16'hCFA0;
defparam \ex_reg_rs1_bypass[11]~48 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[11]~49 (
	.dataa(\ex_reg_rs1_bypass[0]~4_combout ),
	.datab(\ex_reg_rs1_bypass[11]~46_combout ),
	.datac(\ex_reg_rs1_bypass[11]~48_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[11]~49_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[11]~49 .lut_mask = 16'hECEC;
defparam \ex_reg_rs1_bypass[11]~49 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[11]~97 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[11]~q ),
	.datad(\ex_reg_rs1_bypass[11]~49_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[11]~97_combout ),
	.cout());
defparam \alu_io_op1[11]~97 .lut_mask = 16'h6240;
defparam \alu_io_op1[11]~97 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_csr_addr~7 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[31]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_csr_addr~7_combout ),
	.cout());
defparam \ex_csr_addr~7 .lut_mask = 16'h8080;
defparam \ex_csr_addr~7 .sum_lutc_input = "datac";

dffeas \ex_csr_addr[11] (
	.clk(clk_clk),
	.d(\ex_csr_addr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_csr_addr[11]~q ),
	.prn(vcc));
defparam \ex_csr_addr[11] .is_wysiwyg = "true";
defparam \ex_csr_addr[11] .power_up = "low";

cyclone10lp_lcell_comb \_T_3593~0 (
	.dataa(\ex_inst[7]~q ),
	.datab(\ex_ctrl_imm_type.010~q ),
	.datac(\ex_csr_addr[11]~q ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\_T_3593~0_combout ),
	.cout());
defparam \_T_3593~0 .lut_mask = 16'h88B8;
defparam \_T_3593~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_imm_type~21 (
	.dataa(\id_pc[7]~31_combout ),
	.datab(\Equal7~0_combout ),
	.datac(\Equal53~0_combout ),
	.datad(\id_inst[4]~q ),
	.cin(gnd),
	.combout(\ex_ctrl_imm_type~21_combout ),
	.cout());
defparam \ex_ctrl_imm_type~21 .lut_mask = 16'h0040;
defparam \ex_ctrl_imm_type~21 .sum_lutc_input = "datac";

dffeas \ex_ctrl_imm_type.100 (
	.clk(clk_clk),
	.d(\ex_ctrl_imm_type~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_imm_type.100~q ),
	.prn(vcc));
defparam \ex_ctrl_imm_type.100 .is_wysiwyg = "true";
defparam \ex_ctrl_imm_type.100 .power_up = "low";

cyclone10lp_lcell_comb \_T_3593~1 (
	.dataa(\ex_csr_addr[0]~q ),
	.datab(\_T_3593~0_combout ),
	.datac(gnd),
	.datad(\ex_ctrl_imm_type.100~q ),
	.cin(gnd),
	.combout(\_T_3593~1_combout ),
	.cout());
defparam \_T_3593~1 .lut_mask = 16'hAACC;
defparam \_T_3593~1 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a21 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[11]~22_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a21_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_a_first_bit_number = 21;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_b_first_bit_number = 21;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a21 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~11 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a21~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~11_combout ),
	.cout());
defparam \ex_rs_1~11 .lut_mask = 16'h8888;
defparam \ex_rs_1~11 .sum_lutc_input = "datac";

dffeas \ex_rs_1[11] (
	.clk(clk_clk),
	.d(\ex_rs_1~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[11]~q ),
	.prn(vcc));
defparam \ex_rs_1[11] .is_wysiwyg = "true";
defparam \ex_rs_1[11] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[11]~40 (
	.dataa(\ex_reg_rs2_bypass[7]~5_combout ),
	.datab(\ex_rs_1[11]~q ),
	.datac(\ex_reg_rs2_bypass[7]~4_combout ),
	.datad(\wb_alu_out[11]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[11]~40_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[11]~40 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[11]~40 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[11]~41 (
	.dataa(av_readdata_pre_11),
	.datab(\ex_reg_rs2_bypass[7]~5_combout ),
	.datac(\ex_reg_rs2_bypass[11]~40_combout ),
	.datad(\wb_csr_data[11]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[11]~41_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[11]~41 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[11]~41 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[11]~42 (
	.dataa(\mem_alu_out[11]~q ),
	.datab(\ex_reg_rs2_bypass[11]~41_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[11]~42_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[11]~42 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[11]~42 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[11]~50 (
	.dataa(\_T_3681~3_combout ),
	.datab(\mem_csr_data[11]~q ),
	.datac(\ex_reg_rs2_bypass[11]~42_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\alu_io_op2[11]~50_combout ),
	.cout());
defparam \alu_io_op2[11]~50 .lut_mask = 16'hF8F8;
defparam \alu_io_op2[11]~50 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[11]~51 (
	.dataa(\alu_io_op2[5]~43_combout ),
	.datab(\_T_3593~1_combout ),
	.datac(\ex_ctrl_alu_op2.10~q ),
	.datad(\alu_io_op2[11]~50_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[11]~51_combout ),
	.cout());
defparam \alu_io_op2[11]~51 .lut_mask = 16'hA808;
defparam \alu_io_op2[11]~51 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~46 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\alu|_T_123[11]~combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~195_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~46_combout ),
	.cout());
defparam \mem_alu_out~46 .lut_mask = 16'hDAD0;
defparam \mem_alu_out~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~47 (
	.dataa(\alu_io_op1[11]~97_combout ),
	.datab(\alu_io_op2[11]~51_combout ),
	.datac(\mem_alu_out~46_combout ),
	.datad(\alu|LessThan0~0_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~47_combout ),
	.cout());
defparam \mem_alu_out~47 .lut_mask = 16'hF08E;
defparam \mem_alu_out~47 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~48 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[11]~51_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~47_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~48_combout ),
	.cout());
defparam \mem_alu_out~48 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~48 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~49 (
	.dataa(\alu_io_op1[11]~97_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~48_combout ),
	.datad(\alu|ShiftRight0~197_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~49_combout ),
	.cout());
defparam \mem_alu_out~49 .lut_mask = 16'hF838;
defparam \mem_alu_out~49 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~50 (
	.dataa(\mem_alu_out~49_combout ),
	.datab(\alu|_T_3[11]~22_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~50_combout ),
	.cout());
defparam \mem_alu_out~50 .lut_mask = 16'h00AC;
defparam \mem_alu_out~50 .sum_lutc_input = "datac";

dffeas \mem_alu_out[11] (
	.clk(clk_clk),
	.d(\mem_alu_out~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[11]~q ),
	.prn(vcc));
defparam \mem_alu_out[11] .is_wysiwyg = "true";
defparam \mem_alu_out[11] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~9 (
	.dataa(\ex_pc[11]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~9_combout ),
	.cout());
defparam \mem_pc~9 .lut_mask = 16'h8888;
defparam \mem_pc~9 .sum_lutc_input = "datac";

dffeas \mem_pc[11] (
	.clk(clk_clk),
	.d(\mem_pc~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[11]~q ),
	.prn(vcc));
defparam \mem_pc[11] .is_wysiwyg = "true";
defparam \mem_pc[11] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~26 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\_T_3593~1_combout ),
	.datac(\ex_ctrl_imm_type.101~q ),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\mem_imm~26_combout ),
	.cout());
defparam \mem_imm~26 .lut_mask = 16'h0008;
defparam \mem_imm~26 .sum_lutc_input = "datac";

dffeas \mem_imm[11] (
	.clk(clk_clk),
	.d(\mem_imm~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[11]~q ),
	.prn(vcc));
defparam \mem_imm[11] .is_wysiwyg = "true";
defparam \mem_imm[11] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[11]~22 (
	.dataa(\mem_pc[11]~q ),
	.datab(\mem_imm[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[10]~21 ),
	.combout(\_T_3862[11]~22_combout ),
	.cout(\_T_3862[11]~23 ));
defparam \_T_3862[11]~22 .lut_mask = 16'h9617;
defparam \_T_3862[11]~22 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~37 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[11]~22_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[11]~18_combout ),
	.cin(gnd),
	.combout(\pc_cntr~37_combout ),
	.cout());
defparam \pc_cntr~37 .lut_mask = 16'h5E0E;
defparam \pc_cntr~37 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~38 (
	.dataa(\mem_alu_out[11]~q ),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~37_combout ),
	.datad(\csr|mepc[11]~q ),
	.cin(gnd),
	.combout(\pc_cntr~38_combout ),
	.cout());
defparam \pc_cntr~38 .lut_mask = 16'hF838;
defparam \pc_cntr~38 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~39 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~38_combout ),
	.datac(\csr|mtvec[11]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~39_combout ),
	.cout());
defparam \pc_cntr~39 .lut_mask = 16'h88A0;
defparam \pc_cntr~39 .sum_lutc_input = "datac";

dffeas \pc_cntr[11] (
	.clk(clk_clk),
	.d(\pc_cntr~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[11]~q ),
	.prn(vcc));
defparam \pc_cntr[11] .is_wysiwyg = "true";
defparam \pc_cntr[11] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~10 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[11]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~10_combout ),
	.cout());
defparam \id_pc~10 .lut_mask = 16'h8080;
defparam \id_pc~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~10 (
	.dataa(id_pc_12),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~10_combout ),
	.cout());
defparam \ex_pc~10 .lut_mask = 16'h8080;
defparam \ex_pc~10 .sum_lutc_input = "datac";

dffeas \ex_pc[12] (
	.clk(clk_clk),
	.d(\ex_pc~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[12]~q ),
	.prn(vcc));
defparam \ex_pc[12] .is_wysiwyg = "true";
defparam \ex_pc[12] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~10 (
	.dataa(\ex_pc[12]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~10_combout ),
	.cout());
defparam \mem_pc~10 .lut_mask = 16'h8888;
defparam \mem_pc~10 .sum_lutc_input = "datac";

dffeas \mem_pc[12] (
	.clk(clk_clk),
	.d(\mem_pc~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[12]~q ),
	.prn(vcc));
defparam \mem_pc[12] .is_wysiwyg = "true";
defparam \mem_pc[12] .power_up = "low";

cyclone10lp_lcell_comb \ex_inst~11 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[12]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~11_combout ),
	.cout());
defparam \ex_inst~11 .lut_mask = 16'h8080;
defparam \ex_inst~11 .sum_lutc_input = "datac";

dffeas \ex_inst[12] (
	.clk(clk_clk),
	.d(\ex_inst~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[12]~q ),
	.prn(vcc));
defparam \ex_inst[12] .is_wysiwyg = "true";
defparam \ex_inst[12] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~7 (
	.dataa(\ex_csr_addr[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\mem_imm~7_combout ),
	.cout());
defparam \mem_imm~7 .lut_mask = 16'h00AA;
defparam \mem_imm~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb _T_3579(
	.dataa(\ex_ctrl_imm_type.011~q ),
	.datab(\ex_ctrl_imm_type.100~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\_T_3579~combout ),
	.cout());
defparam _T_3579.lut_mask = 16'hEEEE;
defparam _T_3579.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~27 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_inst[12]~q ),
	.datac(\mem_imm~7_combout ),
	.datad(\_T_3579~combout ),
	.cin(gnd),
	.combout(\mem_imm~27_combout ),
	.cout());
defparam \mem_imm~27 .lut_mask = 16'h88A0;
defparam \mem_imm~27 .sum_lutc_input = "datac";

dffeas \mem_imm[12] (
	.clk(clk_clk),
	.d(\mem_imm~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[12]~q ),
	.prn(vcc));
defparam \mem_imm[12] .is_wysiwyg = "true";
defparam \mem_imm[12] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[12]~24 (
	.dataa(\mem_pc[12]~q ),
	.datab(\mem_imm[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[11]~23 ),
	.combout(\_T_3862[12]~24_combout ),
	.cout(\_T_3862[12]~25 ));
defparam \_T_3862[12]~24 .lut_mask = 16'h698E;
defparam \_T_3862[12]~24 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \alu_io_op2[12]~53 (
	.dataa(\ex_inst[12]~q ),
	.datab(\mem_imm~7_combout ),
	.datac(\_T_3579~combout ),
	.datad(\ex_ctrl_alu_op2.10~q ),
	.cin(gnd),
	.combout(\alu_io_op2[12]~53_combout ),
	.cout());
defparam \alu_io_op2[12]~53 .lut_mask = 16'h00AC;
defparam \alu_io_op2[12]~53 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_csr_data~17 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[12]~86_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~17_combout ),
	.cout());
defparam \mem_csr_data~17 .lut_mask = 16'h8888;
defparam \mem_csr_data~17 .sum_lutc_input = "datac";

dffeas \mem_csr_data[12] (
	.clk(clk_clk),
	.d(\mem_csr_data~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[12]~q ),
	.prn(vcc));
defparam \mem_csr_data[12] .is_wysiwyg = "true";
defparam \mem_csr_data[12] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~10 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~10_combout ),
	.cout());
defparam \wb_csr_data~10 .lut_mask = 16'h8888;
defparam \wb_csr_data~10 .sum_lutc_input = "datac";

dffeas \wb_csr_data[12] (
	.clk(clk_clk),
	.d(\wb_csr_data~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[12]~q ),
	.prn(vcc));
defparam \wb_csr_data[12] .is_wysiwyg = "true";
defparam \wb_csr_data[12] .power_up = "low";

cyclone10lp_lcell_comb \npc[12]~20 (
	.dataa(\pc_cntr[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[11]~19 ),
	.combout(\npc[12]~20_combout ),
	.cout(\npc[12]~21 ));
defparam \npc[12]~20 .lut_mask = 16'hA50A;
defparam \npc[12]~20 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~10 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[12]~20_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~10_combout ),
	.cout());
defparam \id_npc~10 .lut_mask = 16'h8080;
defparam \id_npc~10 .sum_lutc_input = "datac";

dffeas \id_npc[12] (
	.clk(clk_clk),
	.d(\id_npc~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[12]~q ),
	.prn(vcc));
defparam \id_npc[12] .is_wysiwyg = "true";
defparam \id_npc[12] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~10 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[12]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~10_combout ),
	.cout());
defparam \ex_npc~10 .lut_mask = 16'h8080;
defparam \ex_npc~10 .sum_lutc_input = "datac";

dffeas \ex_npc[12] (
	.clk(clk_clk),
	.d(\ex_npc~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[12]~q ),
	.prn(vcc));
defparam \ex_npc[12] .is_wysiwyg = "true";
defparam \ex_npc[12] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~8 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~8_combout ),
	.cout());
defparam \mem_npc~8 .lut_mask = 16'h8888;
defparam \mem_npc~8 .sum_lutc_input = "datac";

dffeas \mem_npc[12] (
	.clk(clk_clk),
	.d(\mem_npc~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[12]~q ),
	.prn(vcc));
defparam \mem_npc[12] .is_wysiwyg = "true";
defparam \mem_npc[12] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~8 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~8_combout ),
	.cout());
defparam \wb_npc~8 .lut_mask = 16'h8888;
defparam \wb_npc~8 .sum_lutc_input = "datac";

dffeas \wb_npc[12] (
	.clk(clk_clk),
	.d(\wb_npc~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[12]~q ),
	.prn(vcc));
defparam \wb_npc[12] .is_wysiwyg = "true";
defparam \wb_npc[12] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~10 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~10_combout ),
	.cout());
defparam \wb_alu_out~10 .lut_mask = 16'h8888;
defparam \wb_alu_out~10 .sum_lutc_input = "datac";

dffeas \wb_alu_out[12] (
	.clk(clk_clk),
	.d(\wb_alu_out~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[12]~q ),
	.prn(vcc));
defparam \wb_alu_out[12] .is_wysiwyg = "true";
defparam \wb_alu_out[12] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[12]~23 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[12]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[12]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[12]~23_combout ),
	.cout());
defparam \_T_3543__T_3854_data[12]~23 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[12]~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~61 (
	.dataa(\wb_dmem_read_data[22]~89_combout ),
	.datab(av_readdata_pre_23),
	.datac(\wb_dmem_read_data[22]~90_combout ),
	.datad(\wb_dmem_read_data~60_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~61_combout ),
	.cout());
defparam \wb_dmem_read_data~61 .lut_mask = 16'hE5E0;
defparam \wb_dmem_read_data~61 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~62 (
	.dataa(av_readdata_pre_7),
	.datab(\wb_dmem_read_data[22]~89_combout ),
	.datac(\wb_dmem_read_data~61_combout ),
	.datad(\wb_dmem_read_data~28_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~62_combout ),
	.cout());
defparam \wb_dmem_read_data~62 .lut_mask = 16'hF838;
defparam \wb_dmem_read_data~62 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~63 (
	.dataa(av_readdata_pre_12),
	.datab(\wb_dmem_read_data~62_combout ),
	.datac(\wb_dmem_read_data[14]~45_combout ),
	.datad(\wb_dmem_read_data[14]~47_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~63_combout ),
	.cout());
defparam \wb_dmem_read_data~63 .lut_mask = 16'h00AC;
defparam \wb_dmem_read_data~63 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[12] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[12]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[12] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[12] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[12]~24 (
	.dataa(\wb_csr_data[12]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[12]~23_combout ),
	.datad(\wb_dmem_read_data[12]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[12]~24_combout ),
	.cout());
defparam \_T_3543__T_3854_data[12]~24 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[12]~24 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a20 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[12]~24_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a20_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_a_first_bit_number = 20;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_b_first_bit_number = 20;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a20 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~13 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a20~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~13_combout ),
	.cout());
defparam \ex_rs_1~13 .lut_mask = 16'h8888;
defparam \ex_rs_1~13 .sum_lutc_input = "datac";

dffeas \ex_rs_1[12] (
	.clk(clk_clk),
	.d(\ex_rs_1~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[12]~q ),
	.prn(vcc));
defparam \ex_rs_1[12] .is_wysiwyg = "true";
defparam \ex_rs_1[12] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[12]~47 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_12),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[12]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[12]~47_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[12]~47 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[12]~47 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[12]~48 (
	.dataa(\ex_rs_1[12]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[12]~47_combout ),
	.datad(\wb_csr_data[12]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[12]~48_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[12]~48 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[12]~48 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[12]~49 (
	.dataa(\mem_alu_out[12]~q ),
	.datab(\ex_reg_rs2_bypass[12]~48_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[12]~49_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[12]~49 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[12]~49 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[12]~50 (
	.dataa(\ex_reg_rs2_bypass[12]~49_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[12]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[12]~50_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[12]~50 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[12]~50 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[12]~78 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\alu_io_op2[12]~53_combout ),
	.datad(\ex_reg_rs2_bypass[12]~50_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[12]~78_combout ),
	.cout());
defparam \alu_io_op2[12]~78 .lut_mask = 16'hF8F0;
defparam \alu_io_op2[12]~78 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[12]~50 (
	.dataa(\ex_reg_rs1_bypass[0]~20_combout ),
	.datab(\mem_alu_out[12]~q ),
	.datac(\_T_3634~2_combout ),
	.datad(\mem_csr_data[12]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[12]~50_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[12]~50 .lut_mask = 16'hF888;
defparam \ex_reg_rs1_bypass[12]~50 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a20 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[12]~24_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a20_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_a_first_bit_number = 20;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_b_first_bit_number = 20;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a20 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~12 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a20~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~12_combout ),
	.cout());
defparam \ex_rs_0~12 .lut_mask = 16'h0080;
defparam \ex_rs_0~12 .sum_lutc_input = "datac";

dffeas \ex_rs_0[12] (
	.clk(clk_clk),
	.d(\ex_rs_0~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[12]~q ),
	.prn(vcc));
defparam \ex_rs_0[12] .is_wysiwyg = "true";
defparam \ex_rs_0[12] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[12]~51 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(av_readdata_pre_12),
	.datac(\wb_alu_out[12]~q ),
	.datad(\ex_reg_rs1_bypass[2]~138_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[12]~51_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[12]~51 .lut_mask = 16'hAAD8;
defparam \ex_reg_rs1_bypass[12]~51 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[12]~52 (
	.dataa(\ex_rs_0[12]~q ),
	.datab(\wb_csr_data[12]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\ex_reg_rs1_bypass[12]~51_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[12]~52_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[12]~52 .lut_mask = 16'hCFA0;
defparam \ex_reg_rs1_bypass[12]~52 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[12]~53 (
	.dataa(\ex_reg_rs1_bypass[0]~4_combout ),
	.datab(\ex_reg_rs1_bypass[12]~50_combout ),
	.datac(\ex_reg_rs1_bypass[12]~52_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[12]~53_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[12]~53 .lut_mask = 16'hECEC;
defparam \ex_reg_rs1_bypass[12]~53 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[12]~98 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[12]~q ),
	.datad(\ex_reg_rs1_bypass[12]~53_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[12]~98_combout ),
	.cout());
defparam \alu_io_op1[12]~98 .lut_mask = 16'h6240;
defparam \alu_io_op1[12]~98 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~149 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\alu_io_op2[12]~78_combout ),
	.datad(\alu_io_op1[12]~98_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~149_combout ),
	.cout());
defparam \mem_alu_out~149 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~149 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~150 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~149_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~198_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~150_combout ),
	.cout());
defparam \mem_alu_out~150 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~150 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~51 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[12]~98_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~150_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~51_combout ),
	.cout());
defparam \mem_alu_out~51 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~51 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~52 (
	.dataa(\alu_io_op2[12]~78_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~51_combout ),
	.datad(\alu|ShiftRight0~203_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~52_combout ),
	.cout());
defparam \mem_alu_out~52 .lut_mask = 16'hF838;
defparam \mem_alu_out~52 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~53 (
	.dataa(\mem_alu_out~52_combout ),
	.datab(\alu|_T_3[12]~24_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~53_combout ),
	.cout());
defparam \mem_alu_out~53 .lut_mask = 16'h00AC;
defparam \mem_alu_out~53 .sum_lutc_input = "datac";

dffeas \mem_alu_out[12] (
	.clk(clk_clk),
	.d(\mem_alu_out~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[12]~q ),
	.prn(vcc));
defparam \mem_alu_out[12] .is_wysiwyg = "true";
defparam \mem_alu_out[12] .power_up = "low";

cyclone10lp_lcell_comb \pc_cntr~40 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(\mem_alu_out[12]~q ),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[12]~20_combout ),
	.cin(gnd),
	.combout(\pc_cntr~40_combout ),
	.cout());
defparam \pc_cntr~40 .lut_mask = 16'hDAD0;
defparam \pc_cntr~40 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~41 (
	.dataa(\_T_3862[12]~24_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~40_combout ),
	.datad(\csr|mepc[12]~q ),
	.cin(gnd),
	.combout(\pc_cntr~41_combout ),
	.cout());
defparam \pc_cntr~41 .lut_mask = 16'hF2C2;
defparam \pc_cntr~41 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~42 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~41_combout ),
	.datac(\csr|mtvec[12]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~42_combout ),
	.cout());
defparam \pc_cntr~42 .lut_mask = 16'h88A0;
defparam \pc_cntr~42 .sum_lutc_input = "datac";

dffeas \pc_cntr[12] (
	.clk(clk_clk),
	.d(\pc_cntr~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[12]~q ),
	.prn(vcc));
defparam \pc_cntr[12] .is_wysiwyg = "true";
defparam \pc_cntr[12] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~11 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[12]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~11_combout ),
	.cout());
defparam \id_pc~11 .lut_mask = 16'h8080;
defparam \id_pc~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~11 (
	.dataa(id_pc_13),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~11_combout ),
	.cout());
defparam \ex_pc~11 .lut_mask = 16'h8080;
defparam \ex_pc~11 .sum_lutc_input = "datac";

dffeas \ex_pc[13] (
	.clk(clk_clk),
	.d(\ex_pc~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[13]~q ),
	.prn(vcc));
defparam \ex_pc[13] .is_wysiwyg = "true";
defparam \ex_pc[13] .power_up = "low";

cyclone10lp_lcell_comb \mem_csr_data~18 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[13]~93_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~18_combout ),
	.cout());
defparam \mem_csr_data~18 .lut_mask = 16'h8888;
defparam \mem_csr_data~18 .sum_lutc_input = "datac";

dffeas \mem_csr_data[13] (
	.clk(clk_clk),
	.d(\mem_csr_data~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[13]~q ),
	.prn(vcc));
defparam \mem_csr_data[13] .is_wysiwyg = "true";
defparam \mem_csr_data[13] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[13]~54 (
	.dataa(\ex_reg_rs1_bypass[0]~20_combout ),
	.datab(\mem_alu_out[13]~q ),
	.datac(\_T_3634~2_combout ),
	.datad(\mem_csr_data[13]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[13]~54_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[13]~54 .lut_mask = 16'hF888;
defparam \ex_reg_rs1_bypass[13]~54 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_csr_data~11 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~11_combout ),
	.cout());
defparam \wb_csr_data~11 .lut_mask = 16'h8888;
defparam \wb_csr_data~11 .sum_lutc_input = "datac";

dffeas \wb_csr_data[13] (
	.clk(clk_clk),
	.d(\wb_csr_data~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[13]~q ),
	.prn(vcc));
defparam \wb_csr_data[13] .is_wysiwyg = "true";
defparam \wb_csr_data[13] .power_up = "low";

cyclone10lp_lcell_comb \npc[13]~22 (
	.dataa(\pc_cntr[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[12]~21 ),
	.combout(\npc[13]~22_combout ),
	.cout(\npc[13]~23 ));
defparam \npc[13]~22 .lut_mask = 16'h5A5F;
defparam \npc[13]~22 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~11 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[13]~22_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~11_combout ),
	.cout());
defparam \id_npc~11 .lut_mask = 16'h8080;
defparam \id_npc~11 .sum_lutc_input = "datac";

dffeas \id_npc[13] (
	.clk(clk_clk),
	.d(\id_npc~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[13]~q ),
	.prn(vcc));
defparam \id_npc[13] .is_wysiwyg = "true";
defparam \id_npc[13] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~11 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[13]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~11_combout ),
	.cout());
defparam \ex_npc~11 .lut_mask = 16'h8080;
defparam \ex_npc~11 .sum_lutc_input = "datac";

dffeas \ex_npc[13] (
	.clk(clk_clk),
	.d(\ex_npc~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[13]~q ),
	.prn(vcc));
defparam \ex_npc[13] .is_wysiwyg = "true";
defparam \ex_npc[13] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~9 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~9_combout ),
	.cout());
defparam \mem_npc~9 .lut_mask = 16'h8888;
defparam \mem_npc~9 .sum_lutc_input = "datac";

dffeas \mem_npc[13] (
	.clk(clk_clk),
	.d(\mem_npc~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[13]~q ),
	.prn(vcc));
defparam \mem_npc[13] .is_wysiwyg = "true";
defparam \mem_npc[13] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~9 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~9_combout ),
	.cout());
defparam \wb_npc~9 .lut_mask = 16'h8888;
defparam \wb_npc~9 .sum_lutc_input = "datac";

dffeas \wb_npc[13] (
	.clk(clk_clk),
	.d(\wb_npc~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[13]~q ),
	.prn(vcc));
defparam \wb_npc[13] .is_wysiwyg = "true";
defparam \wb_npc[13] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~11 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~11_combout ),
	.cout());
defparam \wb_alu_out~11 .lut_mask = 16'h8888;
defparam \wb_alu_out~11 .sum_lutc_input = "datac";

dffeas \wb_alu_out[13] (
	.clk(clk_clk),
	.d(\wb_alu_out~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[13]~q ),
	.prn(vcc));
defparam \wb_alu_out[13] .is_wysiwyg = "true";
defparam \wb_alu_out[13] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[13]~25 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[13]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[13]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[13]~25_combout ),
	.cout());
defparam \_T_3543__T_3854_data[13]~25 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[13]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~65 (
	.dataa(\wb_dmem_read_data[22]~90_combout ),
	.datab(av_readdata_pre_7),
	.datac(\wb_dmem_read_data[22]~89_combout ),
	.datad(\wb_dmem_read_data~64_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~65_combout ),
	.cout());
defparam \wb_dmem_read_data~65 .lut_mask = 16'hE5E0;
defparam \wb_dmem_read_data~65 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~66 (
	.dataa(av_readdata_pre_23),
	.datab(\wb_dmem_read_data[22]~90_combout ),
	.datac(\wb_dmem_read_data~65_combout ),
	.datad(\wb_dmem_read_data~28_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~66_combout ),
	.cout());
defparam \wb_dmem_read_data~66 .lut_mask = 16'hF838;
defparam \wb_dmem_read_data~66 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~67 (
	.dataa(av_readdata_pre_13),
	.datab(\wb_dmem_read_data~66_combout ),
	.datac(\wb_dmem_read_data[14]~45_combout ),
	.datad(\wb_dmem_read_data[14]~47_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~67_combout ),
	.cout());
defparam \wb_dmem_read_data~67 .lut_mask = 16'h00AC;
defparam \wb_dmem_read_data~67 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[13] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~67_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[13]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[13] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[13] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[13]~26 (
	.dataa(\wb_npc[13]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[13]~25_combout ),
	.datad(\wb_dmem_read_data[13]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[13]~26_combout ),
	.cout());
defparam \_T_3543__T_3854_data[13]~26 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[13]~26 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a19 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[13]~26_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a19_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_a_first_bit_number = 19;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_b_first_bit_number = 19;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a19 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~13 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a19~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~13_combout ),
	.cout());
defparam \ex_rs_0~13 .lut_mask = 16'h0080;
defparam \ex_rs_0~13 .sum_lutc_input = "datac";

dffeas \ex_rs_0[13] (
	.clk(clk_clk),
	.d(\ex_rs_0~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[13]~q ),
	.prn(vcc));
defparam \ex_rs_0[13] .is_wysiwyg = "true";
defparam \ex_rs_0[13] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[13]~55 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(\ex_rs_0[13]~q ),
	.datac(\wb_alu_out[13]~q ),
	.datad(\ex_reg_rs1_bypass[2]~7_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[13]~55_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[13]~55 .lut_mask = 16'hAAD8;
defparam \ex_reg_rs1_bypass[13]~55 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[13]~56 (
	.dataa(av_readdata_pre_13),
	.datab(\wb_csr_data[13]~q ),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\ex_reg_rs1_bypass[13]~55_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[13]~56_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[13]~56 .lut_mask = 16'hCFA0;
defparam \ex_reg_rs1_bypass[13]~56 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[13]~57 (
	.dataa(\ex_reg_rs1_bypass[0]~4_combout ),
	.datab(\ex_reg_rs1_bypass[13]~54_combout ),
	.datac(\ex_reg_rs1_bypass[13]~56_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[13]~57_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[13]~57 .lut_mask = 16'hECEC;
defparam \ex_reg_rs1_bypass[13]~57 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[13]~99 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[13]~q ),
	.datad(\ex_reg_rs1_bypass[13]~57_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[13]~99_combout ),
	.cout());
defparam \alu_io_op1[13]~99 .lut_mask = 16'h6240;
defparam \alu_io_op1[13]~99 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_inst~10 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[13]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~10_combout ),
	.cout());
defparam \ex_inst~10 .lut_mask = 16'h8080;
defparam \ex_inst~10 .sum_lutc_input = "datac";

dffeas \ex_inst[13] (
	.clk(clk_clk),
	.d(\ex_inst~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[13]~q ),
	.prn(vcc));
defparam \ex_inst[13] .is_wysiwyg = "true";
defparam \ex_inst[13] .power_up = "low";

cyclone10lp_lcell_comb \alu_io_op2[13]~52 (
	.dataa(\ex_inst[13]~q ),
	.datab(\mem_imm~7_combout ),
	.datac(\_T_3579~combout ),
	.datad(\ex_ctrl_alu_op2.10~q ),
	.cin(gnd),
	.combout(\alu_io_op2[13]~52_combout ),
	.cout());
defparam \alu_io_op2[13]~52 .lut_mask = 16'h00AC;
defparam \alu_io_op2[13]~52 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a19 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[13]~26_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a19_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_a_first_bit_number = 19;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_b_first_bit_number = 19;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a19 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~12 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a19~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~12_combout ),
	.cout());
defparam \ex_rs_1~12 .lut_mask = 16'h8888;
defparam \ex_rs_1~12 .sum_lutc_input = "datac";

dffeas \ex_rs_1[13] (
	.clk(clk_clk),
	.d(\ex_rs_1~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[13]~q ),
	.prn(vcc));
defparam \ex_rs_1[13] .is_wysiwyg = "true";
defparam \ex_rs_1[13] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[13]~43 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(\ex_rs_1[13]~q ),
	.datac(\wb_alu_out[13]~q ),
	.datad(\ex_reg_rs2_bypass[7]~5_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[13]~43_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[13]~43 .lut_mask = 16'hAAD8;
defparam \ex_reg_rs2_bypass[13]~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[13]~44 (
	.dataa(av_readdata_pre_13),
	.datab(\wb_csr_data[13]~q ),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\ex_reg_rs2_bypass[13]~43_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[13]~44_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[13]~44 .lut_mask = 16'hCFA0;
defparam \ex_reg_rs2_bypass[13]~44 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[13]~45 (
	.dataa(\mem_alu_out[13]~q ),
	.datab(\_T_3686~0_combout ),
	.datac(\_T_3681~3_combout ),
	.datad(\ex_reg_rs2_bypass[13]~44_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[13]~45_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[13]~45 .lut_mask = 16'h0B08;
defparam \ex_reg_rs2_bypass[13]~45 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[13]~46 (
	.dataa(\ex_reg_rs2_bypass[13]~45_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[13]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[13]~46_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[13]~46 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[13]~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[13]~77 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\alu_io_op2[13]~52_combout ),
	.datad(\ex_reg_rs2_bypass[13]~46_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[13]~77_combout ),
	.cout());
defparam \alu_io_op2[13]~77 .lut_mask = 16'hF8F0;
defparam \alu_io_op2[13]~77 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~54 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\alu|_T_123[13]~combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~249_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~54_combout ),
	.cout());
defparam \mem_alu_out~54 .lut_mask = 16'hDAD0;
defparam \mem_alu_out~54 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~55 (
	.dataa(\alu_io_op1[13]~99_combout ),
	.datab(\alu_io_op2[13]~77_combout ),
	.datac(\mem_alu_out~54_combout ),
	.datad(\alu|LessThan0~0_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~55_combout ),
	.cout());
defparam \mem_alu_out~55 .lut_mask = 16'hF08E;
defparam \mem_alu_out~55 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~56 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[13]~77_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~55_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~56_combout ),
	.cout());
defparam \mem_alu_out~56 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~56 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~57 (
	.dataa(\alu_io_op1[13]~99_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~56_combout ),
	.datad(\alu|ShiftRight0~209_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~57_combout ),
	.cout());
defparam \mem_alu_out~57 .lut_mask = 16'hF838;
defparam \mem_alu_out~57 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~58 (
	.dataa(\mem_alu_out~57_combout ),
	.datab(\alu|_T_3[13]~26_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~58_combout ),
	.cout());
defparam \mem_alu_out~58 .lut_mask = 16'h00AC;
defparam \mem_alu_out~58 .sum_lutc_input = "datac";

dffeas \mem_alu_out[13] (
	.clk(clk_clk),
	.d(\mem_alu_out~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[13]~q ),
	.prn(vcc));
defparam \mem_alu_out[13] .is_wysiwyg = "true";
defparam \mem_alu_out[13] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~11 (
	.dataa(\ex_pc[13]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~11_combout ),
	.cout());
defparam \mem_pc~11 .lut_mask = 16'h8888;
defparam \mem_pc~11 .sum_lutc_input = "datac";

dffeas \mem_pc[13] (
	.clk(clk_clk),
	.d(\mem_pc~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[13]~q ),
	.prn(vcc));
defparam \mem_pc[13] .is_wysiwyg = "true";
defparam \mem_pc[13] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~28 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_inst[13]~q ),
	.datac(\mem_imm~7_combout ),
	.datad(\_T_3579~combout ),
	.cin(gnd),
	.combout(\mem_imm~28_combout ),
	.cout());
defparam \mem_imm~28 .lut_mask = 16'h88A0;
defparam \mem_imm~28 .sum_lutc_input = "datac";

dffeas \mem_imm[13] (
	.clk(clk_clk),
	.d(\mem_imm~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[13]~q ),
	.prn(vcc));
defparam \mem_imm[13] .is_wysiwyg = "true";
defparam \mem_imm[13] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[13]~26 (
	.dataa(\mem_pc[13]~q ),
	.datab(\mem_imm[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[12]~25 ),
	.combout(\_T_3862[13]~26_combout ),
	.cout(\_T_3862[13]~27 ));
defparam \_T_3862[13]~26 .lut_mask = 16'h9617;
defparam \_T_3862[13]~26 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~43 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[13]~26_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[13]~22_combout ),
	.cin(gnd),
	.combout(\pc_cntr~43_combout ),
	.cout());
defparam \pc_cntr~43 .lut_mask = 16'h5E0E;
defparam \pc_cntr~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~44 (
	.dataa(\mem_alu_out[13]~q ),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~43_combout ),
	.datad(\csr|mepc[13]~q ),
	.cin(gnd),
	.combout(\pc_cntr~44_combout ),
	.cout());
defparam \pc_cntr~44 .lut_mask = 16'hF838;
defparam \pc_cntr~44 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~45 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~44_combout ),
	.datac(\csr|mtvec[13]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~45_combout ),
	.cout());
defparam \pc_cntr~45 .lut_mask = 16'h88A0;
defparam \pc_cntr~45 .sum_lutc_input = "datac";

dffeas \pc_cntr[13] (
	.clk(clk_clk),
	.d(\pc_cntr~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[13]~q ),
	.prn(vcc));
defparam \pc_cntr[13] .is_wysiwyg = "true";
defparam \pc_cntr[13] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~12 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[13]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~12_combout ),
	.cout());
defparam \id_pc~12 .lut_mask = 16'h8080;
defparam \id_pc~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~12 (
	.dataa(id_pc_14),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~12_combout ),
	.cout());
defparam \ex_pc~12 .lut_mask = 16'h8080;
defparam \ex_pc~12 .sum_lutc_input = "datac";

dffeas \ex_pc[14] (
	.clk(clk_clk),
	.d(\ex_pc~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[14]~q ),
	.prn(vcc));
defparam \ex_pc[14] .is_wysiwyg = "true";
defparam \ex_pc[14] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~12 (
	.dataa(\ex_pc[14]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~12_combout ),
	.cout());
defparam \mem_pc~12 .lut_mask = 16'h8888;
defparam \mem_pc~12 .sum_lutc_input = "datac";

dffeas \mem_pc[14] (
	.clk(clk_clk),
	.d(\mem_pc~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[14]~q ),
	.prn(vcc));
defparam \mem_pc[14] .is_wysiwyg = "true";
defparam \mem_pc[14] .power_up = "low";

cyclone10lp_lcell_comb \ex_inst~12 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_inst[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_inst~12_combout ),
	.cout());
defparam \ex_inst~12 .lut_mask = 16'h8080;
defparam \ex_inst~12 .sum_lutc_input = "datac";

dffeas \ex_inst[14] (
	.clk(clk_clk),
	.d(\ex_inst~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_inst[14]~q ),
	.prn(vcc));
defparam \ex_inst[14] .is_wysiwyg = "true";
defparam \ex_inst[14] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~29 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_inst[14]~q ),
	.datac(\mem_imm~7_combout ),
	.datad(\_T_3579~combout ),
	.cin(gnd),
	.combout(\mem_imm~29_combout ),
	.cout());
defparam \mem_imm~29 .lut_mask = 16'h88A0;
defparam \mem_imm~29 .sum_lutc_input = "datac";

dffeas \mem_imm[14] (
	.clk(clk_clk),
	.d(\mem_imm~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[14]~q ),
	.prn(vcc));
defparam \mem_imm[14] .is_wysiwyg = "true";
defparam \mem_imm[14] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[14]~28 (
	.dataa(\mem_pc[14]~q ),
	.datab(\mem_imm[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[13]~27 ),
	.combout(\_T_3862[14]~28_combout ),
	.cout(\_T_3862[14]~29 ));
defparam \_T_3862[14]~28 .lut_mask = 16'h698E;
defparam \_T_3862[14]~28 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \alu_io_op2[14]~54 (
	.dataa(\ex_inst[14]~q ),
	.datab(\mem_imm~7_combout ),
	.datac(\_T_3579~combout ),
	.datad(\ex_ctrl_alu_op2.10~q ),
	.cin(gnd),
	.combout(\alu_io_op2[14]~54_combout ),
	.cout());
defparam \alu_io_op2[14]~54 .lut_mask = 16'h00AC;
defparam \alu_io_op2[14]~54 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_csr_data~19 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[14]~100_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~19_combout ),
	.cout());
defparam \mem_csr_data~19 .lut_mask = 16'h8888;
defparam \mem_csr_data~19 .sum_lutc_input = "datac";

dffeas \mem_csr_data[14] (
	.clk(clk_clk),
	.d(\mem_csr_data~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[14]~q ),
	.prn(vcc));
defparam \mem_csr_data[14] .is_wysiwyg = "true";
defparam \mem_csr_data[14] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~12 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~12_combout ),
	.cout());
defparam \wb_csr_data~12 .lut_mask = 16'h8888;
defparam \wb_csr_data~12 .sum_lutc_input = "datac";

dffeas \wb_csr_data[14] (
	.clk(clk_clk),
	.d(\wb_csr_data~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[14]~q ),
	.prn(vcc));
defparam \wb_csr_data[14] .is_wysiwyg = "true";
defparam \wb_csr_data[14] .power_up = "low";

cyclone10lp_lcell_comb \npc[14]~24 (
	.dataa(\pc_cntr[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[13]~23 ),
	.combout(\npc[14]~24_combout ),
	.cout(\npc[14]~25 ));
defparam \npc[14]~24 .lut_mask = 16'hA50A;
defparam \npc[14]~24 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~12 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[14]~24_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~12_combout ),
	.cout());
defparam \id_npc~12 .lut_mask = 16'h8080;
defparam \id_npc~12 .sum_lutc_input = "datac";

dffeas \id_npc[14] (
	.clk(clk_clk),
	.d(\id_npc~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[14]~q ),
	.prn(vcc));
defparam \id_npc[14] .is_wysiwyg = "true";
defparam \id_npc[14] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~12 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~12_combout ),
	.cout());
defparam \ex_npc~12 .lut_mask = 16'h8080;
defparam \ex_npc~12 .sum_lutc_input = "datac";

dffeas \ex_npc[14] (
	.clk(clk_clk),
	.d(\ex_npc~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[14]~q ),
	.prn(vcc));
defparam \ex_npc[14] .is_wysiwyg = "true";
defparam \ex_npc[14] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~10 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~10_combout ),
	.cout());
defparam \mem_npc~10 .lut_mask = 16'h8888;
defparam \mem_npc~10 .sum_lutc_input = "datac";

dffeas \mem_npc[14] (
	.clk(clk_clk),
	.d(\mem_npc~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[14]~q ),
	.prn(vcc));
defparam \mem_npc[14] .is_wysiwyg = "true";
defparam \mem_npc[14] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~10 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~10_combout ),
	.cout());
defparam \wb_npc~10 .lut_mask = 16'h8888;
defparam \wb_npc~10 .sum_lutc_input = "datac";

dffeas \wb_npc[14] (
	.clk(clk_clk),
	.d(\wb_npc~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[14]~q ),
	.prn(vcc));
defparam \wb_npc[14] .is_wysiwyg = "true";
defparam \wb_npc[14] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~12 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~12_combout ),
	.cout());
defparam \wb_alu_out~12 .lut_mask = 16'h8888;
defparam \wb_alu_out~12 .sum_lutc_input = "datac";

dffeas \wb_alu_out[14] (
	.clk(clk_clk),
	.d(\wb_alu_out~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[14]~q ),
	.prn(vcc));
defparam \wb_alu_out[14] .is_wysiwyg = "true";
defparam \wb_alu_out[14] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[14]~27 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[14]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[14]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[14]~27_combout ),
	.cout());
defparam \_T_3543__T_3854_data[14]~27 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[14]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~69 (
	.dataa(\wb_dmem_read_data[22]~89_combout ),
	.datab(av_readdata_pre_23),
	.datac(\wb_dmem_read_data[22]~90_combout ),
	.datad(\wb_dmem_read_data~68_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~69_combout ),
	.cout());
defparam \wb_dmem_read_data~69 .lut_mask = 16'hE5E0;
defparam \wb_dmem_read_data~69 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~70 (
	.dataa(av_readdata_pre_7),
	.datab(\wb_dmem_read_data[22]~89_combout ),
	.datac(\wb_dmem_read_data~69_combout ),
	.datad(\wb_dmem_read_data~28_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~70_combout ),
	.cout());
defparam \wb_dmem_read_data~70 .lut_mask = 16'hF838;
defparam \wb_dmem_read_data~70 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~71 (
	.dataa(av_readdata_pre_14),
	.datab(\wb_dmem_read_data~70_combout ),
	.datac(\wb_dmem_read_data[14]~45_combout ),
	.datad(\wb_dmem_read_data[14]~47_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~71_combout ),
	.cout());
defparam \wb_dmem_read_data~71 .lut_mask = 16'h00AC;
defparam \wb_dmem_read_data~71 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[14] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~71_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[14]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[14] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[14] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[14]~28 (
	.dataa(\wb_csr_data[14]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[14]~27_combout ),
	.datad(\wb_dmem_read_data[14]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[14]~28_combout ),
	.cout());
defparam \_T_3543__T_3854_data[14]~28 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[14]~28 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a18 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[14]~28_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a18_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_a_first_bit_number = 18;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_b_first_bit_number = 18;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a18 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~14 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a18~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~14_combout ),
	.cout());
defparam \ex_rs_1~14 .lut_mask = 16'h8888;
defparam \ex_rs_1~14 .sum_lutc_input = "datac";

dffeas \ex_rs_1[14] (
	.clk(clk_clk),
	.d(\ex_rs_1~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[14]~q ),
	.prn(vcc));
defparam \ex_rs_1[14] .is_wysiwyg = "true";
defparam \ex_rs_1[14] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[14]~51 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_14),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[14]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[14]~51_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[14]~51 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[14]~51 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[14]~52 (
	.dataa(\ex_rs_1[14]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[14]~51_combout ),
	.datad(\wb_csr_data[14]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[14]~52_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[14]~52 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[14]~52 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[14]~53 (
	.dataa(\mem_alu_out[14]~q ),
	.datab(\ex_reg_rs2_bypass[14]~52_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[14]~53_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[14]~53 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[14]~53 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[14]~54 (
	.dataa(\ex_reg_rs2_bypass[14]~53_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[14]~54_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[14]~54 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[14]~54 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[14]~79 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\alu_io_op2[14]~54_combout ),
	.datad(\ex_reg_rs2_bypass[14]~54_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[14]~79_combout ),
	.cout());
defparam \alu_io_op2[14]~79 .lut_mask = 16'hF8F0;
defparam \alu_io_op2[14]~79 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[14]~58 (
	.dataa(\ex_reg_rs1_bypass[0]~20_combout ),
	.datab(\mem_alu_out[14]~q ),
	.datac(\_T_3634~2_combout ),
	.datad(\mem_csr_data[14]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[14]~58_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[14]~58 .lut_mask = 16'hF888;
defparam \ex_reg_rs1_bypass[14]~58 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a18 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[14]~28_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a18_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_a_first_bit_number = 18;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_b_first_bit_number = 18;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a18 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~14 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a18~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~14_combout ),
	.cout());
defparam \ex_rs_0~14 .lut_mask = 16'h0080;
defparam \ex_rs_0~14 .sum_lutc_input = "datac";

dffeas \ex_rs_0[14] (
	.clk(clk_clk),
	.d(\ex_rs_0~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[14]~q ),
	.prn(vcc));
defparam \ex_rs_0[14] .is_wysiwyg = "true";
defparam \ex_rs_0[14] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[14]~59 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(av_readdata_pre_14),
	.datac(\wb_alu_out[14]~q ),
	.datad(\ex_reg_rs1_bypass[2]~138_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[14]~59_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[14]~59 .lut_mask = 16'hAAD8;
defparam \ex_reg_rs1_bypass[14]~59 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[14]~60 (
	.dataa(\ex_rs_0[14]~q ),
	.datab(\wb_csr_data[14]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\ex_reg_rs1_bypass[14]~59_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[14]~60_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[14]~60 .lut_mask = 16'hCFA0;
defparam \ex_reg_rs1_bypass[14]~60 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[14]~61 (
	.dataa(\ex_reg_rs1_bypass[0]~4_combout ),
	.datab(\ex_reg_rs1_bypass[14]~58_combout ),
	.datac(\ex_reg_rs1_bypass[14]~60_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[14]~61_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[14]~61 .lut_mask = 16'hECEC;
defparam \ex_reg_rs1_bypass[14]~61 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[14]~100 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[14]~q ),
	.datad(\ex_reg_rs1_bypass[14]~61_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[14]~100_combout ),
	.cout());
defparam \alu_io_op1[14]~100 .lut_mask = 16'h6240;
defparam \alu_io_op1[14]~100 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~147 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\alu_io_op2[14]~79_combout ),
	.datad(\alu_io_op1[14]~100_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~147_combout ),
	.cout());
defparam \mem_alu_out~147 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~147 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~148 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~147_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~250_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~148_combout ),
	.cout());
defparam \mem_alu_out~148 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~148 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~59 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[14]~100_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~148_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~59_combout ),
	.cout());
defparam \mem_alu_out~59 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~59 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~60 (
	.dataa(\alu_io_op2[14]~79_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~59_combout ),
	.datad(\alu|ShiftRight0~216_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~60_combout ),
	.cout());
defparam \mem_alu_out~60 .lut_mask = 16'hF838;
defparam \mem_alu_out~60 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~61 (
	.dataa(\mem_alu_out~60_combout ),
	.datab(\alu|_T_3[14]~28_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~61_combout ),
	.cout());
defparam \mem_alu_out~61 .lut_mask = 16'h00AC;
defparam \mem_alu_out~61 .sum_lutc_input = "datac";

dffeas \mem_alu_out[14] (
	.clk(clk_clk),
	.d(\mem_alu_out~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[14]~q ),
	.prn(vcc));
defparam \mem_alu_out[14] .is_wysiwyg = "true";
defparam \mem_alu_out[14] .power_up = "low";

cyclone10lp_lcell_comb \pc_cntr~46 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(\mem_alu_out[14]~q ),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[14]~24_combout ),
	.cin(gnd),
	.combout(\pc_cntr~46_combout ),
	.cout());
defparam \pc_cntr~46 .lut_mask = 16'hDAD0;
defparam \pc_cntr~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~47 (
	.dataa(\_T_3862[14]~28_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~46_combout ),
	.datad(\csr|mepc[14]~q ),
	.cin(gnd),
	.combout(\pc_cntr~47_combout ),
	.cout());
defparam \pc_cntr~47 .lut_mask = 16'hF2C2;
defparam \pc_cntr~47 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~48 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~47_combout ),
	.datac(\csr|mtvec[14]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~48_combout ),
	.cout());
defparam \pc_cntr~48 .lut_mask = 16'h88A0;
defparam \pc_cntr~48 .sum_lutc_input = "datac";

dffeas \pc_cntr[14] (
	.clk(clk_clk),
	.d(\pc_cntr~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[14]~q ),
	.prn(vcc));
defparam \pc_cntr[14] .is_wysiwyg = "true";
defparam \pc_cntr[14] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~13 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~13_combout ),
	.cout());
defparam \id_pc~13 .lut_mask = 16'h8080;
defparam \id_pc~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~13 (
	.dataa(id_pc_15),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~13_combout ),
	.cout());
defparam \ex_pc~13 .lut_mask = 16'h8080;
defparam \ex_pc~13 .sum_lutc_input = "datac";

dffeas \ex_pc[15] (
	.clk(clk_clk),
	.d(\ex_pc~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[15]~q ),
	.prn(vcc));
defparam \ex_pc[15] .is_wysiwyg = "true";
defparam \ex_pc[15] .power_up = "low";

cyclone10lp_lcell_comb \mem_csr_data~20 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[15]~107_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~20_combout ),
	.cout());
defparam \mem_csr_data~20 .lut_mask = 16'h8888;
defparam \mem_csr_data~20 .sum_lutc_input = "datac";

dffeas \mem_csr_data[15] (
	.clk(clk_clk),
	.d(\mem_csr_data~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[15]~q ),
	.prn(vcc));
defparam \mem_csr_data[15] .is_wysiwyg = "true";
defparam \mem_csr_data[15] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[15]~62 (
	.dataa(\ex_reg_rs1_bypass[0]~20_combout ),
	.datab(\mem_alu_out[15]~q ),
	.datac(\_T_3634~2_combout ),
	.datad(\mem_csr_data[15]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[15]~62_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[15]~62 .lut_mask = 16'hF888;
defparam \ex_reg_rs1_bypass[15]~62 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_csr_data~13 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~13_combout ),
	.cout());
defparam \wb_csr_data~13 .lut_mask = 16'h8888;
defparam \wb_csr_data~13 .sum_lutc_input = "datac";

dffeas \wb_csr_data[15] (
	.clk(clk_clk),
	.d(\wb_csr_data~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[15]~q ),
	.prn(vcc));
defparam \wb_csr_data[15] .is_wysiwyg = "true";
defparam \wb_csr_data[15] .power_up = "low";

cyclone10lp_lcell_comb \npc[15]~26 (
	.dataa(\pc_cntr[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[14]~25 ),
	.combout(\npc[15]~26_combout ),
	.cout(\npc[15]~27 ));
defparam \npc[15]~26 .lut_mask = 16'h5A5F;
defparam \npc[15]~26 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~13 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[15]~26_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~13_combout ),
	.cout());
defparam \id_npc~13 .lut_mask = 16'h8080;
defparam \id_npc~13 .sum_lutc_input = "datac";

dffeas \id_npc[15] (
	.clk(clk_clk),
	.d(\id_npc~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[15]~q ),
	.prn(vcc));
defparam \id_npc[15] .is_wysiwyg = "true";
defparam \id_npc[15] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~13 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[15]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~13_combout ),
	.cout());
defparam \ex_npc~13 .lut_mask = 16'h8080;
defparam \ex_npc~13 .sum_lutc_input = "datac";

dffeas \ex_npc[15] (
	.clk(clk_clk),
	.d(\ex_npc~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[15]~q ),
	.prn(vcc));
defparam \ex_npc[15] .is_wysiwyg = "true";
defparam \ex_npc[15] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~11 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~11_combout ),
	.cout());
defparam \mem_npc~11 .lut_mask = 16'h8888;
defparam \mem_npc~11 .sum_lutc_input = "datac";

dffeas \mem_npc[15] (
	.clk(clk_clk),
	.d(\mem_npc~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[15]~q ),
	.prn(vcc));
defparam \mem_npc[15] .is_wysiwyg = "true";
defparam \mem_npc[15] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~11 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~11_combout ),
	.cout());
defparam \wb_npc~11 .lut_mask = 16'h8888;
defparam \wb_npc~11 .sum_lutc_input = "datac";

dffeas \wb_npc[15] (
	.clk(clk_clk),
	.d(\wb_npc~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[15]~q ),
	.prn(vcc));
defparam \wb_npc[15] .is_wysiwyg = "true";
defparam \wb_npc[15] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~13 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~13_combout ),
	.cout());
defparam \wb_alu_out~13 .lut_mask = 16'h8888;
defparam \wb_alu_out~13 .sum_lutc_input = "datac";

dffeas \wb_alu_out[15] (
	.clk(clk_clk),
	.d(\wb_alu_out~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[15]~q ),
	.prn(vcc));
defparam \wb_alu_out[15] .is_wysiwyg = "true";
defparam \wb_alu_out[15] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[15]~29 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[15]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[15]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[15]~29_combout ),
	.cout());
defparam \_T_3543__T_3854_data[15]~29 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[15]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~72 (
	.dataa(av_readdata_pre_15),
	.datab(\mem_ctrl_mask_type[0]~q ),
	.datac(\mem_ctrl_mask_type[1]~q ),
	.datad(mem_ctrl_mem_wr01),
	.cin(gnd),
	.combout(\wb_dmem_read_data~72_combout ),
	.cout());
defparam \wb_dmem_read_data~72 .lut_mask = 16'h82AA;
defparam \wb_dmem_read_data~72 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~91 (
	.dataa(mem_alu_out_0),
	.datab(mem_alu_out_1),
	.datac(\wb_dmem_read_data~28_combout ),
	.datad(av_readdata_pre_23),
	.cin(gnd),
	.combout(\wb_dmem_read_data~91_combout ),
	.cout());
defparam \wb_dmem_read_data~91 .lut_mask = 16'hE4A0;
defparam \wb_dmem_read_data~91 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal69~0 (
	.dataa(mem_alu_out_0),
	.datab(mem_alu_out_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal69~0_combout ),
	.cout());
defparam \Equal69~0 .lut_mask = 16'hEEEE;
defparam \Equal69~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~39 (
	.dataa(Equal68),
	.datab(\wb_dmem_read_data~91_combout ),
	.datac(av_readdata_pre_7),
	.datad(\Equal69~0_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~39_combout ),
	.cout());
defparam \wb_dmem_read_data~39 .lut_mask = 16'h88A8;
defparam \wb_dmem_read_data~39 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~73 (
	.dataa(\mem_ctrl_mask_type[1]~q ),
	.datab(\wb_dmem_read_data~28_combout ),
	.datac(mem_alu_out_0),
	.datad(\mem_ctrl_mask_type[0]~q ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~73_combout ),
	.cout());
defparam \wb_dmem_read_data~73 .lut_mask = 16'h0008;
defparam \wb_dmem_read_data~73 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~74 (
	.dataa(\wb_dmem_read_data~72_combout ),
	.datab(mem_ctrl_mem_wr01),
	.datac(\wb_dmem_read_data~39_combout ),
	.datad(\wb_dmem_read_data~73_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~74_combout ),
	.cout());
defparam \wb_dmem_read_data~74 .lut_mask = 16'hEEEA;
defparam \wb_dmem_read_data~74 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[15] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[15]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[15] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[15] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[15]~30 (
	.dataa(\wb_npc[15]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[15]~29_combout ),
	.datad(\wb_dmem_read_data[15]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[15]~30_combout ),
	.cout());
defparam \_T_3543__T_3854_data[15]~30 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[15]~30 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a17 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[15]~30_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a17_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_a_first_bit_number = 17;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_b_first_bit_number = 17;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a17 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~15 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a17~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~15_combout ),
	.cout());
defparam \ex_rs_0~15 .lut_mask = 16'h0080;
defparam \ex_rs_0~15 .sum_lutc_input = "datac";

dffeas \ex_rs_0[15] (
	.clk(clk_clk),
	.d(\ex_rs_0~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[15]~q ),
	.prn(vcc));
defparam \ex_rs_0[15] .is_wysiwyg = "true";
defparam \ex_rs_0[15] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[15]~63 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(\ex_rs_0[15]~q ),
	.datac(\wb_alu_out[15]~q ),
	.datad(\ex_reg_rs1_bypass[2]~7_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[15]~63_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[15]~63 .lut_mask = 16'hAAD8;
defparam \ex_reg_rs1_bypass[15]~63 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[15]~64 (
	.dataa(av_readdata_pre_15),
	.datab(\wb_csr_data[15]~q ),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\ex_reg_rs1_bypass[15]~63_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[15]~64_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[15]~64 .lut_mask = 16'hCFA0;
defparam \ex_reg_rs1_bypass[15]~64 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[15]~65 (
	.dataa(\ex_reg_rs1_bypass[0]~4_combout ),
	.datab(\ex_reg_rs1_bypass[15]~62_combout ),
	.datac(\ex_reg_rs1_bypass[15]~64_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[15]~65_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[15]~65 .lut_mask = 16'hECEC;
defparam \ex_reg_rs1_bypass[15]~65 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[15]~101 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[15]~q ),
	.datad(\ex_reg_rs1_bypass[15]~65_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[15]~101_combout ),
	.cout());
defparam \alu_io_op1[15]~101 .lut_mask = 16'h6240;
defparam \alu_io_op1[15]~101 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[15]~55 (
	.dataa(\ex_inst[15]~q ),
	.datab(\mem_imm~7_combout ),
	.datac(\_T_3579~combout ),
	.datad(\ex_ctrl_alu_op2.10~q ),
	.cin(gnd),
	.combout(\alu_io_op2[15]~55_combout ),
	.cout());
defparam \alu_io_op2[15]~55 .lut_mask = 16'h00AC;
defparam \alu_io_op2[15]~55 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a17 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[15]~30_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a17_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_a_first_bit_number = 17;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_b_first_bit_number = 17;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a17 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~15 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a17~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~15_combout ),
	.cout());
defparam \ex_rs_1~15 .lut_mask = 16'h8888;
defparam \ex_rs_1~15 .sum_lutc_input = "datac";

dffeas \ex_rs_1[15] (
	.clk(clk_clk),
	.d(\ex_rs_1~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[15]~q ),
	.prn(vcc));
defparam \ex_rs_1[15] .is_wysiwyg = "true";
defparam \ex_rs_1[15] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[15]~55 (
	.dataa(\ex_reg_rs2_bypass[7]~5_combout ),
	.datab(\ex_rs_1[15]~q ),
	.datac(\ex_reg_rs2_bypass[7]~4_combout ),
	.datad(\wb_alu_out[15]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[15]~55_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[15]~55 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[15]~55 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[15]~56 (
	.dataa(av_readdata_pre_15),
	.datab(\ex_reg_rs2_bypass[7]~5_combout ),
	.datac(\ex_reg_rs2_bypass[15]~55_combout ),
	.datad(\wb_csr_data[15]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[15]~56_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[15]~56 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[15]~56 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[15]~57 (
	.dataa(\mem_alu_out[15]~q ),
	.datab(\ex_reg_rs2_bypass[15]~56_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[15]~57_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[15]~57 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[15]~57 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[15]~58 (
	.dataa(\ex_reg_rs2_bypass[15]~57_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[15]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[15]~58_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[15]~58 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[15]~58 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[15]~92 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\alu_io_op2[15]~55_combout ),
	.datad(\ex_reg_rs2_bypass[15]~58_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[15]~92_combout ),
	.cout());
defparam \alu_io_op2[15]~92 .lut_mask = 16'hF8F0;
defparam \alu_io_op2[15]~92 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~62 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\alu|_T_123[15]~combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~217_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~62_combout ),
	.cout());
defparam \mem_alu_out~62 .lut_mask = 16'hDAD0;
defparam \mem_alu_out~62 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~63 (
	.dataa(\alu_io_op1[15]~101_combout ),
	.datab(\alu_io_op2[15]~92_combout ),
	.datac(\mem_alu_out~62_combout ),
	.datad(\alu|LessThan0~0_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~63_combout ),
	.cout());
defparam \mem_alu_out~63 .lut_mask = 16'hF08E;
defparam \mem_alu_out~63 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~64 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[15]~92_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~63_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~64_combout ),
	.cout());
defparam \mem_alu_out~64 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~64 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~65 (
	.dataa(\alu_io_op1[15]~101_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~64_combout ),
	.datad(\alu|ShiftRight0~222_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~65_combout ),
	.cout());
defparam \mem_alu_out~65 .lut_mask = 16'hF838;
defparam \mem_alu_out~65 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~66 (
	.dataa(\mem_alu_out~65_combout ),
	.datab(\alu|_T_3[15]~30_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~66_combout ),
	.cout());
defparam \mem_alu_out~66 .lut_mask = 16'h00AC;
defparam \mem_alu_out~66 .sum_lutc_input = "datac";

dffeas \mem_alu_out[15] (
	.clk(clk_clk),
	.d(\mem_alu_out~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[15]~q ),
	.prn(vcc));
defparam \mem_alu_out[15] .is_wysiwyg = "true";
defparam \mem_alu_out[15] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~13 (
	.dataa(\ex_pc[15]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~13_combout ),
	.cout());
defparam \mem_pc~13 .lut_mask = 16'h8888;
defparam \mem_pc~13 .sum_lutc_input = "datac";

dffeas \mem_pc[15] (
	.clk(clk_clk),
	.d(\mem_pc~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[15]~q ),
	.prn(vcc));
defparam \mem_pc[15] .is_wysiwyg = "true";
defparam \mem_pc[15] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~30 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_inst[15]~q ),
	.datac(\mem_imm~7_combout ),
	.datad(\_T_3579~combout ),
	.cin(gnd),
	.combout(\mem_imm~30_combout ),
	.cout());
defparam \mem_imm~30 .lut_mask = 16'h88A0;
defparam \mem_imm~30 .sum_lutc_input = "datac";

dffeas \mem_imm[15] (
	.clk(clk_clk),
	.d(\mem_imm~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[15]~q ),
	.prn(vcc));
defparam \mem_imm[15] .is_wysiwyg = "true";
defparam \mem_imm[15] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[15]~30 (
	.dataa(\mem_pc[15]~q ),
	.datab(\mem_imm[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[14]~29 ),
	.combout(\_T_3862[15]~30_combout ),
	.cout(\_T_3862[15]~31 ));
defparam \_T_3862[15]~30 .lut_mask = 16'h9617;
defparam \_T_3862[15]~30 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~49 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[15]~30_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[15]~26_combout ),
	.cin(gnd),
	.combout(\pc_cntr~49_combout ),
	.cout());
defparam \pc_cntr~49 .lut_mask = 16'h5E0E;
defparam \pc_cntr~49 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~50 (
	.dataa(\mem_alu_out[15]~q ),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~49_combout ),
	.datad(\csr|mepc[15]~q ),
	.cin(gnd),
	.combout(\pc_cntr~50_combout ),
	.cout());
defparam \pc_cntr~50 .lut_mask = 16'hF838;
defparam \pc_cntr~50 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~51 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~50_combout ),
	.datac(\csr|mtvec[15]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~51_combout ),
	.cout());
defparam \pc_cntr~51 .lut_mask = 16'h88A0;
defparam \pc_cntr~51 .sum_lutc_input = "datac";

dffeas \pc_cntr[15] (
	.clk(clk_clk),
	.d(\pc_cntr~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[15]~q ),
	.prn(vcc));
defparam \pc_cntr[15] .is_wysiwyg = "true";
defparam \pc_cntr[15] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~14 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[15]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~14_combout ),
	.cout());
defparam \id_pc~14 .lut_mask = 16'h8080;
defparam \id_pc~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~14 (
	.dataa(id_pc_16),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~14_combout ),
	.cout());
defparam \ex_pc~14 .lut_mask = 16'h8080;
defparam \ex_pc~14 .sum_lutc_input = "datac";

dffeas \ex_pc[16] (
	.clk(clk_clk),
	.d(\ex_pc~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[16]~q ),
	.prn(vcc));
defparam \ex_pc[16] .is_wysiwyg = "true";
defparam \ex_pc[16] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~14 (
	.dataa(\ex_pc[16]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~14_combout ),
	.cout());
defparam \mem_pc~14 .lut_mask = 16'h8888;
defparam \mem_pc~14 .sum_lutc_input = "datac";

dffeas \mem_pc[16] (
	.clk(clk_clk),
	.d(\mem_pc~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[16]~q ),
	.prn(vcc));
defparam \mem_pc[16] .is_wysiwyg = "true";
defparam \mem_pc[16] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~31 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_inst[16]~q ),
	.datac(\mem_imm~7_combout ),
	.datad(\_T_3579~combout ),
	.cin(gnd),
	.combout(\mem_imm~31_combout ),
	.cout());
defparam \mem_imm~31 .lut_mask = 16'h88A0;
defparam \mem_imm~31 .sum_lutc_input = "datac";

dffeas \mem_imm[16] (
	.clk(clk_clk),
	.d(\mem_imm~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[16]~q ),
	.prn(vcc));
defparam \mem_imm[16] .is_wysiwyg = "true";
defparam \mem_imm[16] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[16]~32 (
	.dataa(\mem_pc[16]~q ),
	.datab(\mem_imm[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[15]~31 ),
	.combout(\_T_3862[16]~32_combout ),
	.cout(\_T_3862[16]~33 ));
defparam \_T_3862[16]~32 .lut_mask = 16'h698E;
defparam \_T_3862[16]~32 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \alu_io_op2[16]~57 (
	.dataa(\ex_inst[16]~q ),
	.datab(\mem_imm~7_combout ),
	.datac(\_T_3579~combout ),
	.datad(\ex_ctrl_alu_op2.10~q ),
	.cin(gnd),
	.combout(\alu_io_op2[16]~57_combout ),
	.cout());
defparam \alu_io_op2[16]~57 .lut_mask = 16'h00AC;
defparam \alu_io_op2[16]~57 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_csr_data~21 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[16]~114_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~21_combout ),
	.cout());
defparam \mem_csr_data~21 .lut_mask = 16'h8888;
defparam \mem_csr_data~21 .sum_lutc_input = "datac";

dffeas \mem_csr_data[16] (
	.clk(clk_clk),
	.d(\mem_csr_data~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[16]~q ),
	.prn(vcc));
defparam \mem_csr_data[16] .is_wysiwyg = "true";
defparam \mem_csr_data[16] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~14 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~14_combout ),
	.cout());
defparam \wb_csr_data~14 .lut_mask = 16'h8888;
defparam \wb_csr_data~14 .sum_lutc_input = "datac";

dffeas \wb_csr_data[16] (
	.clk(clk_clk),
	.d(\wb_csr_data~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[16]~q ),
	.prn(vcc));
defparam \wb_csr_data[16] .is_wysiwyg = "true";
defparam \wb_csr_data[16] .power_up = "low";

cyclone10lp_lcell_comb \npc[16]~28 (
	.dataa(\pc_cntr[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[15]~27 ),
	.combout(\npc[16]~28_combout ),
	.cout(\npc[16]~29 ));
defparam \npc[16]~28 .lut_mask = 16'hA50A;
defparam \npc[16]~28 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~14 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[16]~28_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~14_combout ),
	.cout());
defparam \id_npc~14 .lut_mask = 16'h8080;
defparam \id_npc~14 .sum_lutc_input = "datac";

dffeas \id_npc[16] (
	.clk(clk_clk),
	.d(\id_npc~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[16]~q ),
	.prn(vcc));
defparam \id_npc[16] .is_wysiwyg = "true";
defparam \id_npc[16] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~14 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[16]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~14_combout ),
	.cout());
defparam \ex_npc~14 .lut_mask = 16'h8080;
defparam \ex_npc~14 .sum_lutc_input = "datac";

dffeas \ex_npc[16] (
	.clk(clk_clk),
	.d(\ex_npc~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[16]~q ),
	.prn(vcc));
defparam \ex_npc[16] .is_wysiwyg = "true";
defparam \ex_npc[16] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~12 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~12_combout ),
	.cout());
defparam \mem_npc~12 .lut_mask = 16'h8888;
defparam \mem_npc~12 .sum_lutc_input = "datac";

dffeas \mem_npc[16] (
	.clk(clk_clk),
	.d(\mem_npc~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[16]~q ),
	.prn(vcc));
defparam \mem_npc[16] .is_wysiwyg = "true";
defparam \mem_npc[16] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~12 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~12_combout ),
	.cout());
defparam \wb_npc~12 .lut_mask = 16'h8888;
defparam \wb_npc~12 .sum_lutc_input = "datac";

dffeas \wb_npc[16] (
	.clk(clk_clk),
	.d(\wb_npc~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[16]~q ),
	.prn(vcc));
defparam \wb_npc[16] .is_wysiwyg = "true";
defparam \wb_npc[16] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~14 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~14_combout ),
	.cout());
defparam \wb_alu_out~14 .lut_mask = 16'h8888;
defparam \wb_alu_out~14 .sum_lutc_input = "datac";

dffeas \wb_alu_out[16] (
	.clk(clk_clk),
	.d(\wb_alu_out~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[16]~q ),
	.prn(vcc));
defparam \wb_alu_out[16] .is_wysiwyg = "true";
defparam \wb_alu_out[16] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[16]~31 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[16]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[16]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[16]~31_combout ),
	.cout());
defparam \_T_3543__T_3854_data[16]~31 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[16]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~23 (
	.dataa(mem_ctrl_mem_wr01),
	.datab(gnd),
	.datac(\mem_ctrl_mask_type[0]~q ),
	.datad(\mem_ctrl_mask_type[1]~q ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~23_combout ),
	.cout());
defparam \wb_dmem_read_data~23 .lut_mask = 16'h0AA0;
defparam \wb_dmem_read_data~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_wb_sel~20 (
	.dataa(\id_inst[5]~q ),
	.datab(\id_inst[6]~q ),
	.datac(\ex_ctrl_mask_type~1_combout ),
	.datad(\Equal9~1_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_wb_sel~20_combout ),
	.cout());
defparam \ex_ctrl_wb_sel~20 .lut_mask = 16'hE0F0;
defparam \ex_ctrl_wb_sel~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mask_type~7 (
	.dataa(\ex_ctrl_wb_sel~20_combout ),
	.datab(\ex_ctrl_mask_type~0_combout ),
	.datac(\_GEN_15~2_combout ),
	.datad(\ex_ctrl_mask_type~2_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_mask_type~7_combout ),
	.cout());
defparam \ex_ctrl_mask_type~7 .lut_mask = 16'h0080;
defparam \ex_ctrl_mask_type~7 .sum_lutc_input = "datac";

dffeas \ex_ctrl_mask_type[2] (
	.clk(clk_clk),
	.d(\ex_ctrl_mask_type~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_mask_type[2]~q ),
	.prn(vcc));
defparam \ex_ctrl_mask_type[2] .is_wysiwyg = "true";
defparam \ex_ctrl_mask_type[2] .power_up = "low";

cyclone10lp_lcell_comb \mem_ctrl_mask_type~1 (
	.dataa(\ex_ctrl_mask_type[2]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_ctrl_mask_type~1_combout ),
	.cout());
defparam \mem_ctrl_mask_type~1 .lut_mask = 16'h8888;
defparam \mem_ctrl_mask_type~1 .sum_lutc_input = "datac";

dffeas \mem_ctrl_mask_type[2] (
	.clk(clk_clk),
	.d(\mem_ctrl_mask_type~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_ctrl_mask_type[2]~q ),
	.prn(vcc));
defparam \mem_ctrl_mask_type[2] .is_wysiwyg = "true";
defparam \mem_ctrl_mask_type[2] .power_up = "low";

cyclone10lp_lcell_comb \wb_dmem_read_data[22]~24 (
	.dataa(\mem_ctrl_mask_type[1]~q ),
	.datab(mem_alu_out_0),
	.datac(\mem_ctrl_mask_type[2]~q ),
	.datad(\mem_ctrl_mask_type[0]~q ),
	.cin(gnd),
	.combout(\wb_dmem_read_data[22]~24_combout ),
	.cout());
defparam \wb_dmem_read_data[22]~24 .lut_mask = 16'h0002;
defparam \wb_dmem_read_data[22]~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[22]~25 (
	.dataa(\Equal69~0_combout ),
	.datab(\mem_ctrl_mask_type[1]~q ),
	.datac(\mem_ctrl_mask_type[2]~q ),
	.datad(\mem_ctrl_mask_type[0]~q ),
	.cin(gnd),
	.combout(\wb_dmem_read_data[22]~25_combout ),
	.cout());
defparam \wb_dmem_read_data[22]~25 .lut_mask = 16'h0008;
defparam \wb_dmem_read_data[22]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~26 (
	.dataa(\wb_dmem_read_data[22]~24_combout ),
	.datab(av_readdata_pre_31),
	.datac(av_readdata_pre_15),
	.datad(\wb_dmem_read_data[22]~25_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~26_combout ),
	.cout());
defparam \wb_dmem_read_data~26 .lut_mask = 16'h88A0;
defparam \wb_dmem_read_data~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~34 (
	.dataa(\wb_dmem_read_data[22]~90_combout ),
	.datab(av_readdata_pre_7),
	.datac(\wb_dmem_read_data[22]~89_combout ),
	.datad(\wb_dmem_read_data~26_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~34_combout ),
	.cout());
defparam \wb_dmem_read_data~34 .lut_mask = 16'hE5E0;
defparam \wb_dmem_read_data~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~35 (
	.dataa(av_readdata_pre_23),
	.datab(\wb_dmem_read_data[22]~90_combout ),
	.datac(\wb_dmem_read_data~34_combout ),
	.datad(\wb_dmem_read_data~28_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~35_combout ),
	.cout());
defparam \wb_dmem_read_data~35 .lut_mask = 16'hF838;
defparam \wb_dmem_read_data~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal68~1 (
	.dataa(\mem_ctrl_mask_type[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_ctrl_mask_type[1]~q ),
	.cin(gnd),
	.combout(\Equal68~1_combout ),
	.cout());
defparam \Equal68~1 .lut_mask = 16'h00AA;
defparam \Equal68~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~36 (
	.dataa(\wb_dmem_read_data~23_combout ),
	.datab(\wb_dmem_read_data~35_combout ),
	.datac(\mem_ctrl_mask_type[2]~q ),
	.datad(\Equal68~1_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~36_combout ),
	.cout());
defparam \wb_dmem_read_data~36 .lut_mask = 16'h0888;
defparam \wb_dmem_read_data~36 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[22]~31 (
	.dataa(\mem_ctrl_mask_type[2]~q ),
	.datab(\mem_ctrl_mask_type[0]~q ),
	.datac(mem_ctrl_mem_wr01),
	.datad(\mem_ctrl_mask_type[1]~q ),
	.cin(gnd),
	.combout(\wb_dmem_read_data[22]~31_combout ),
	.cout());
defparam \wb_dmem_read_data[22]~31 .lut_mask = 16'h0080;
defparam \wb_dmem_read_data[22]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[22]~32 (
	.dataa(\wb_dmem_read_data[22]~31_combout ),
	.datab(mem_alu_out_0),
	.datac(mem_alu_out_1),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\wb_dmem_read_data[22]~32_combout ),
	.cout());
defparam \wb_dmem_read_data[22]~32 .lut_mask = 16'h2AFF;
defparam \wb_dmem_read_data[22]~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~75 (
	.dataa(\wb_dmem_read_data~36_combout ),
	.datab(av_readdata_pre_16),
	.datac(\wb_dmem_read_data~23_combout ),
	.datad(\wb_dmem_read_data[22]~32_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~75_combout ),
	.cout());
defparam \wb_dmem_read_data~75 .lut_mask = 16'h00AE;
defparam \wb_dmem_read_data~75 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[16] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~75_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[16]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[16] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[16] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[16]~32 (
	.dataa(\wb_csr_data[16]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[16]~31_combout ),
	.datad(\wb_dmem_read_data[16]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[16]~32_combout ),
	.cout());
defparam \_T_3543__T_3854_data[16]~32 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[16]~32 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a16 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[16]~32_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a16_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_a_first_bit_number = 16;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_b_first_bit_number = 16;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a16 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~17 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a16~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~17_combout ),
	.cout());
defparam \ex_rs_1~17 .lut_mask = 16'h8888;
defparam \ex_rs_1~17 .sum_lutc_input = "datac";

dffeas \ex_rs_1[16] (
	.clk(clk_clk),
	.d(\ex_rs_1~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[16]~q ),
	.prn(vcc));
defparam \ex_rs_1[16] .is_wysiwyg = "true";
defparam \ex_rs_1[16] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[16]~63 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_16),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[16]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[16]~63_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[16]~63 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[16]~63 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[16]~64 (
	.dataa(\ex_rs_1[16]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[16]~63_combout ),
	.datad(\wb_csr_data[16]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[16]~64_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[16]~64 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[16]~64 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[16]~65 (
	.dataa(\mem_alu_out[16]~q ),
	.datab(\ex_reg_rs2_bypass[16]~64_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[16]~65_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[16]~65 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[16]~65 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[16]~66 (
	.dataa(\ex_reg_rs2_bypass[16]~65_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[16]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[16]~66_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[16]~66 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[16]~66 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[16]~81 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\alu_io_op2[16]~57_combout ),
	.datad(\ex_reg_rs2_bypass[16]~66_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[16]~81_combout ),
	.cout());
defparam \alu_io_op2[16]~81 .lut_mask = 16'hF8F0;
defparam \alu_io_op2[16]~81 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[16]~66 (
	.dataa(\ex_reg_rs1_bypass[0]~20_combout ),
	.datab(\mem_alu_out[16]~q ),
	.datac(\_T_3634~2_combout ),
	.datad(\mem_csr_data[16]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[16]~66_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[16]~66 .lut_mask = 16'hF888;
defparam \ex_reg_rs1_bypass[16]~66 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a16 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[16]~32_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a16_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_a_first_bit_number = 16;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_b_first_bit_number = 16;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a16 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~16 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a16~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~16_combout ),
	.cout());
defparam \ex_rs_0~16 .lut_mask = 16'h0080;
defparam \ex_rs_0~16 .sum_lutc_input = "datac";

dffeas \ex_rs_0[16] (
	.clk(clk_clk),
	.d(\ex_rs_0~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[16]~q ),
	.prn(vcc));
defparam \ex_rs_0[16] .is_wysiwyg = "true";
defparam \ex_rs_0[16] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[16]~67 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(av_readdata_pre_16),
	.datac(\wb_alu_out[16]~q ),
	.datad(\ex_reg_rs1_bypass[2]~138_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[16]~67_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[16]~67 .lut_mask = 16'hAAD8;
defparam \ex_reg_rs1_bypass[16]~67 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[16]~68 (
	.dataa(\ex_rs_0[16]~q ),
	.datab(\wb_csr_data[16]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\ex_reg_rs1_bypass[16]~67_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[16]~68_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[16]~68 .lut_mask = 16'hCFA0;
defparam \ex_reg_rs1_bypass[16]~68 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[16]~69 (
	.dataa(\ex_reg_rs1_bypass[0]~4_combout ),
	.datab(\ex_reg_rs1_bypass[16]~66_combout ),
	.datac(\ex_reg_rs1_bypass[16]~68_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[16]~69_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[16]~69 .lut_mask = 16'hECEC;
defparam \ex_reg_rs1_bypass[16]~69 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[16]~102 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[16]~q ),
	.datad(\ex_reg_rs1_bypass[16]~69_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[16]~102_combout ),
	.cout());
defparam \alu_io_op1[16]~102 .lut_mask = 16'h6240;
defparam \alu_io_op1[16]~102 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~145 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\alu_io_op2[16]~81_combout ),
	.datad(\alu_io_op1[16]~102_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~145_combout ),
	.cout());
defparam \mem_alu_out~145 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~145 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~146 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~145_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~222_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~146_combout ),
	.cout());
defparam \mem_alu_out~146 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~146 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~67 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[16]~102_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~146_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~67_combout ),
	.cout());
defparam \mem_alu_out~67 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~67 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~68 (
	.dataa(\alu_io_op2[16]~81_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~67_combout ),
	.datad(\alu|ShiftRight0~217_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~68_combout ),
	.cout());
defparam \mem_alu_out~68 .lut_mask = 16'hF838;
defparam \mem_alu_out~68 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~69 (
	.dataa(\mem_alu_out~68_combout ),
	.datab(\alu|_T_3[16]~32_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~69_combout ),
	.cout());
defparam \mem_alu_out~69 .lut_mask = 16'h00AC;
defparam \mem_alu_out~69 .sum_lutc_input = "datac";

dffeas \mem_alu_out[16] (
	.clk(clk_clk),
	.d(\mem_alu_out~69_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[16]~q ),
	.prn(vcc));
defparam \mem_alu_out[16] .is_wysiwyg = "true";
defparam \mem_alu_out[16] .power_up = "low";

cyclone10lp_lcell_comb \pc_cntr~52 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(\mem_alu_out[16]~q ),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[16]~28_combout ),
	.cin(gnd),
	.combout(\pc_cntr~52_combout ),
	.cout());
defparam \pc_cntr~52 .lut_mask = 16'hDAD0;
defparam \pc_cntr~52 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~53 (
	.dataa(\_T_3862[16]~32_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~52_combout ),
	.datad(\csr|mepc[16]~q ),
	.cin(gnd),
	.combout(\pc_cntr~53_combout ),
	.cout());
defparam \pc_cntr~53 .lut_mask = 16'hF2C2;
defparam \pc_cntr~53 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~54 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~53_combout ),
	.datac(\csr|mtvec[16]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~54_combout ),
	.cout());
defparam \pc_cntr~54 .lut_mask = 16'h88A0;
defparam \pc_cntr~54 .sum_lutc_input = "datac";

dffeas \pc_cntr[16] (
	.clk(clk_clk),
	.d(\pc_cntr~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[16]~q ),
	.prn(vcc));
defparam \pc_cntr[16] .is_wysiwyg = "true";
defparam \pc_cntr[16] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~15 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[16]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~15_combout ),
	.cout());
defparam \id_pc~15 .lut_mask = 16'h8080;
defparam \id_pc~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~15 (
	.dataa(id_pc_17),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~15_combout ),
	.cout());
defparam \ex_pc~15 .lut_mask = 16'h8080;
defparam \ex_pc~15 .sum_lutc_input = "datac";

dffeas \ex_pc[17] (
	.clk(clk_clk),
	.d(\ex_pc~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[17]~q ),
	.prn(vcc));
defparam \ex_pc[17] .is_wysiwyg = "true";
defparam \ex_pc[17] .power_up = "low";

cyclone10lp_lcell_comb \npc[17]~30 (
	.dataa(\pc_cntr[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[16]~29 ),
	.combout(\npc[17]~30_combout ),
	.cout(\npc[17]~31 ));
defparam \npc[17]~30 .lut_mask = 16'h5A5F;
defparam \npc[17]~30 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~15 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[17]~30_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~15_combout ),
	.cout());
defparam \id_npc~15 .lut_mask = 16'h8080;
defparam \id_npc~15 .sum_lutc_input = "datac";

dffeas \id_npc[17] (
	.clk(clk_clk),
	.d(\id_npc~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[17]~q ),
	.prn(vcc));
defparam \id_npc[17] .is_wysiwyg = "true";
defparam \id_npc[17] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~15 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[17]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~15_combout ),
	.cout());
defparam \ex_npc~15 .lut_mask = 16'h8080;
defparam \ex_npc~15 .sum_lutc_input = "datac";

dffeas \ex_npc[17] (
	.clk(clk_clk),
	.d(\ex_npc~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[17]~q ),
	.prn(vcc));
defparam \ex_npc[17] .is_wysiwyg = "true";
defparam \ex_npc[17] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~13 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~13_combout ),
	.cout());
defparam \mem_npc~13 .lut_mask = 16'h8888;
defparam \mem_npc~13 .sum_lutc_input = "datac";

dffeas \mem_npc[17] (
	.clk(clk_clk),
	.d(\mem_npc~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[17]~q ),
	.prn(vcc));
defparam \mem_npc[17] .is_wysiwyg = "true";
defparam \mem_npc[17] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~13 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~13_combout ),
	.cout());
defparam \wb_npc~13 .lut_mask = 16'h8888;
defparam \wb_npc~13 .sum_lutc_input = "datac";

dffeas \wb_npc[17] (
	.clk(clk_clk),
	.d(\wb_npc~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[17]~q ),
	.prn(vcc));
defparam \wb_npc[17] .is_wysiwyg = "true";
defparam \wb_npc[17] .power_up = "low";

cyclone10lp_lcell_comb \mem_csr_data~22 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[17]~121_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~22_combout ),
	.cout());
defparam \mem_csr_data~22 .lut_mask = 16'h8888;
defparam \mem_csr_data~22 .sum_lutc_input = "datac";

dffeas \mem_csr_data[17] (
	.clk(clk_clk),
	.d(\mem_csr_data~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[17]~q ),
	.prn(vcc));
defparam \mem_csr_data[17] .is_wysiwyg = "true";
defparam \mem_csr_data[17] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~15 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~15_combout ),
	.cout());
defparam \wb_csr_data~15 .lut_mask = 16'h8888;
defparam \wb_csr_data~15 .sum_lutc_input = "datac";

dffeas \wb_csr_data[17] (
	.clk(clk_clk),
	.d(\wb_csr_data~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[17]~q ),
	.prn(vcc));
defparam \wb_csr_data[17] .is_wysiwyg = "true";
defparam \wb_csr_data[17] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~15 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~15_combout ),
	.cout());
defparam \wb_alu_out~15 .lut_mask = 16'h8888;
defparam \wb_alu_out~15 .sum_lutc_input = "datac";

dffeas \wb_alu_out[17] (
	.clk(clk_clk),
	.d(\wb_alu_out~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[17]~q ),
	.prn(vcc));
defparam \wb_alu_out[17] .is_wysiwyg = "true";
defparam \wb_alu_out[17] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[17]~33 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[17]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[17]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[17]~33_combout ),
	.cout());
defparam \_T_3543__T_3854_data[17]~33 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[17]~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~27 (
	.dataa(\wb_dmem_read_data[22]~89_combout ),
	.datab(av_readdata_pre_23),
	.datac(\wb_dmem_read_data[22]~90_combout ),
	.datad(\wb_dmem_read_data~26_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~27_combout ),
	.cout());
defparam \wb_dmem_read_data~27 .lut_mask = 16'hE5E0;
defparam \wb_dmem_read_data~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~29 (
	.dataa(av_readdata_pre_7),
	.datab(\wb_dmem_read_data[22]~89_combout ),
	.datac(\wb_dmem_read_data~27_combout ),
	.datad(\wb_dmem_read_data~28_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~29_combout ),
	.cout());
defparam \wb_dmem_read_data~29 .lut_mask = 16'hF838;
defparam \wb_dmem_read_data~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~30 (
	.dataa(\wb_dmem_read_data~23_combout ),
	.datab(\wb_dmem_read_data~29_combout ),
	.datac(\mem_ctrl_mask_type[2]~q ),
	.datad(\Equal68~1_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~30_combout ),
	.cout());
defparam \wb_dmem_read_data~30 .lut_mask = 16'h0888;
defparam \wb_dmem_read_data~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~76 (
	.dataa(\wb_dmem_read_data~30_combout ),
	.datab(av_readdata_pre_17),
	.datac(\wb_dmem_read_data~23_combout ),
	.datad(\wb_dmem_read_data[22]~32_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~76_combout ),
	.cout());
defparam \wb_dmem_read_data~76 .lut_mask = 16'h00AE;
defparam \wb_dmem_read_data~76 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[17] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[17]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[17] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[17] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[17]~34 (
	.dataa(\wb_npc[17]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[17]~33_combout ),
	.datad(\wb_dmem_read_data[17]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[17]~34_combout ),
	.cout());
defparam \_T_3543__T_3854_data[17]~34 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[17]~34 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a15 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[17]~34_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a15_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_a_first_bit_number = 15;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_b_first_bit_number = 15;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a15 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~17 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a15~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~17_combout ),
	.cout());
defparam \ex_rs_0~17 .lut_mask = 16'h0080;
defparam \ex_rs_0~17 .sum_lutc_input = "datac";

dffeas \ex_rs_0[17] (
	.clk(clk_clk),
	.d(\ex_rs_0~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[17]~q ),
	.prn(vcc));
defparam \ex_rs_0[17] .is_wysiwyg = "true";
defparam \ex_rs_0[17] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[17]~70 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(\ex_rs_0[17]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\wb_alu_out[17]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[17]~70_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[17]~70 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[17]~70 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[17]~71 (
	.dataa(av_readdata_pre_17),
	.datab(\ex_reg_rs1_bypass[2]~7_combout ),
	.datac(\ex_reg_rs1_bypass[17]~70_combout ),
	.datad(\wb_csr_data[17]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[17]~71_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[17]~71 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[17]~71 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[17]~72 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[17]~71_combout ),
	.datad(\mem_csr_data[17]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[17]~72_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[17]~72 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[17]~72 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[17]~73 (
	.dataa(\ex_reg_rs1_bypass[17]~72_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[17]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[17]~73_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[17]~73 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[17]~73 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[17]~103 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[17]~q ),
	.datad(\ex_reg_rs1_bypass[17]~73_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[17]~103_combout ),
	.cout());
defparam \alu_io_op1[17]~103 .lut_mask = 16'h6240;
defparam \alu_io_op1[17]~103 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[17]~56 (
	.dataa(\ex_inst[17]~q ),
	.datab(\mem_imm~7_combout ),
	.datac(\_T_3579~combout ),
	.datad(\ex_ctrl_alu_op2.10~q ),
	.cin(gnd),
	.combout(\alu_io_op2[17]~56_combout ),
	.cout());
defparam \alu_io_op2[17]~56 .lut_mask = 16'h00AC;
defparam \alu_io_op2[17]~56 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a15 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[17]~34_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_a_first_bit_number = 15;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_b_first_bit_number = 15;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a15 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~16 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a15~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~16_combout ),
	.cout());
defparam \ex_rs_1~16 .lut_mask = 16'h8888;
defparam \ex_rs_1~16 .sum_lutc_input = "datac";

dffeas \ex_rs_1[17] (
	.clk(clk_clk),
	.d(\ex_rs_1~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[17]~q ),
	.prn(vcc));
defparam \ex_rs_1[17] .is_wysiwyg = "true";
defparam \ex_rs_1[17] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[17]~59 (
	.dataa(\ex_reg_rs2_bypass[7]~5_combout ),
	.datab(\ex_rs_1[17]~q ),
	.datac(\ex_reg_rs2_bypass[7]~4_combout ),
	.datad(\wb_alu_out[17]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[17]~59_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[17]~59 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[17]~59 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[17]~60 (
	.dataa(av_readdata_pre_17),
	.datab(\ex_reg_rs2_bypass[7]~5_combout ),
	.datac(\ex_reg_rs2_bypass[17]~59_combout ),
	.datad(\wb_csr_data[17]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[17]~60_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[17]~60 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[17]~60 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[17]~61 (
	.dataa(\mem_alu_out[17]~q ),
	.datab(\ex_reg_rs2_bypass[17]~60_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[17]~61_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[17]~61 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[17]~61 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[17]~62 (
	.dataa(\ex_reg_rs2_bypass[17]~61_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[17]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[17]~62_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[17]~62 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[17]~62 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[17]~80 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\alu_io_op2[17]~56_combout ),
	.datad(\ex_reg_rs2_bypass[17]~62_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[17]~80_combout ),
	.cout());
defparam \alu_io_op2[17]~80 .lut_mask = 16'hF8F0;
defparam \alu_io_op2[17]~80 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~70 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\alu|_T_123[17]~combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~216_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~70_combout ),
	.cout());
defparam \mem_alu_out~70 .lut_mask = 16'hDAD0;
defparam \mem_alu_out~70 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~71 (
	.dataa(\alu_io_op1[17]~103_combout ),
	.datab(\alu_io_op2[17]~80_combout ),
	.datac(\mem_alu_out~70_combout ),
	.datad(\alu|LessThan0~0_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~71_combout ),
	.cout());
defparam \mem_alu_out~71 .lut_mask = 16'hF08E;
defparam \mem_alu_out~71 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~72 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[17]~80_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~71_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~72_combout ),
	.cout());
defparam \mem_alu_out~72 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~72 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~73 (
	.dataa(\alu_io_op1[17]~103_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~72_combout ),
	.datad(\alu|ShiftRight0~250_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~73_combout ),
	.cout());
defparam \mem_alu_out~73 .lut_mask = 16'hF838;
defparam \mem_alu_out~73 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~74 (
	.dataa(\mem_alu_out~73_combout ),
	.datab(\alu|_T_3[17]~34_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~74_combout ),
	.cout());
defparam \mem_alu_out~74 .lut_mask = 16'h00AC;
defparam \mem_alu_out~74 .sum_lutc_input = "datac";

dffeas \mem_alu_out[17] (
	.clk(clk_clk),
	.d(\mem_alu_out~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[17]~q ),
	.prn(vcc));
defparam \mem_alu_out[17] .is_wysiwyg = "true";
defparam \mem_alu_out[17] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~15 (
	.dataa(\ex_pc[17]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~15_combout ),
	.cout());
defparam \mem_pc~15 .lut_mask = 16'h8888;
defparam \mem_pc~15 .sum_lutc_input = "datac";

dffeas \mem_pc[17] (
	.clk(clk_clk),
	.d(\mem_pc~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[17]~q ),
	.prn(vcc));
defparam \mem_pc[17] .is_wysiwyg = "true";
defparam \mem_pc[17] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~32 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_inst[17]~q ),
	.datac(\mem_imm~7_combout ),
	.datad(\_T_3579~combout ),
	.cin(gnd),
	.combout(\mem_imm~32_combout ),
	.cout());
defparam \mem_imm~32 .lut_mask = 16'h88A0;
defparam \mem_imm~32 .sum_lutc_input = "datac";

dffeas \mem_imm[17] (
	.clk(clk_clk),
	.d(\mem_imm~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[17]~q ),
	.prn(vcc));
defparam \mem_imm[17] .is_wysiwyg = "true";
defparam \mem_imm[17] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[17]~34 (
	.dataa(\mem_pc[17]~q ),
	.datab(\mem_imm[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[16]~33 ),
	.combout(\_T_3862[17]~34_combout ),
	.cout(\_T_3862[17]~35 ));
defparam \_T_3862[17]~34 .lut_mask = 16'h9617;
defparam \_T_3862[17]~34 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~55 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[17]~34_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[17]~30_combout ),
	.cin(gnd),
	.combout(\pc_cntr~55_combout ),
	.cout());
defparam \pc_cntr~55 .lut_mask = 16'h5E0E;
defparam \pc_cntr~55 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~56 (
	.dataa(\mem_alu_out[17]~q ),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~55_combout ),
	.datad(\csr|mepc[17]~q ),
	.cin(gnd),
	.combout(\pc_cntr~56_combout ),
	.cout());
defparam \pc_cntr~56 .lut_mask = 16'hF838;
defparam \pc_cntr~56 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~57 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~56_combout ),
	.datac(\csr|mtvec[17]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~57_combout ),
	.cout());
defparam \pc_cntr~57 .lut_mask = 16'h88A0;
defparam \pc_cntr~57 .sum_lutc_input = "datac";

dffeas \pc_cntr[17] (
	.clk(clk_clk),
	.d(\pc_cntr~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[17]~q ),
	.prn(vcc));
defparam \pc_cntr[17] .is_wysiwyg = "true";
defparam \pc_cntr[17] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~16 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[17]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~16_combout ),
	.cout());
defparam \id_pc~16 .lut_mask = 16'h8080;
defparam \id_pc~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~16 (
	.dataa(id_pc_18),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~16_combout ),
	.cout());
defparam \ex_pc~16 .lut_mask = 16'h8080;
defparam \ex_pc~16 .sum_lutc_input = "datac";

dffeas \ex_pc[18] (
	.clk(clk_clk),
	.d(\ex_pc~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[18]~q ),
	.prn(vcc));
defparam \ex_pc[18] .is_wysiwyg = "true";
defparam \ex_pc[18] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~16 (
	.dataa(\ex_pc[18]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~16_combout ),
	.cout());
defparam \mem_pc~16 .lut_mask = 16'h8888;
defparam \mem_pc~16 .sum_lutc_input = "datac";

dffeas \mem_pc[18] (
	.clk(clk_clk),
	.d(\mem_pc~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[18]~q ),
	.prn(vcc));
defparam \mem_pc[18] .is_wysiwyg = "true";
defparam \mem_pc[18] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~33 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_inst[18]~q ),
	.datac(\mem_imm~7_combout ),
	.datad(\_T_3579~combout ),
	.cin(gnd),
	.combout(\mem_imm~33_combout ),
	.cout());
defparam \mem_imm~33 .lut_mask = 16'h88A0;
defparam \mem_imm~33 .sum_lutc_input = "datac";

dffeas \mem_imm[18] (
	.clk(clk_clk),
	.d(\mem_imm~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[18]~q ),
	.prn(vcc));
defparam \mem_imm[18] .is_wysiwyg = "true";
defparam \mem_imm[18] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[18]~36 (
	.dataa(\mem_pc[18]~q ),
	.datab(\mem_imm[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[17]~35 ),
	.combout(\_T_3862[18]~36_combout ),
	.cout(\_T_3862[18]~37 ));
defparam \_T_3862[18]~36 .lut_mask = 16'h698E;
defparam \_T_3862[18]~36 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \alu_io_op2[18]~58 (
	.dataa(\ex_inst[18]~q ),
	.datab(\mem_imm~7_combout ),
	.datac(\_T_3579~combout ),
	.datad(\ex_ctrl_alu_op2.10~q ),
	.cin(gnd),
	.combout(\alu_io_op2[18]~58_combout ),
	.cout());
defparam \alu_io_op2[18]~58 .lut_mask = 16'h00AC;
defparam \alu_io_op2[18]~58 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_csr_data~23 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[18]~128_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~23_combout ),
	.cout());
defparam \mem_csr_data~23 .lut_mask = 16'h8888;
defparam \mem_csr_data~23 .sum_lutc_input = "datac";

dffeas \mem_csr_data[18] (
	.clk(clk_clk),
	.d(\mem_csr_data~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[18]~q ),
	.prn(vcc));
defparam \mem_csr_data[18] .is_wysiwyg = "true";
defparam \mem_csr_data[18] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~16 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~16_combout ),
	.cout());
defparam \wb_csr_data~16 .lut_mask = 16'h8888;
defparam \wb_csr_data~16 .sum_lutc_input = "datac";

dffeas \wb_csr_data[18] (
	.clk(clk_clk),
	.d(\wb_csr_data~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[18]~q ),
	.prn(vcc));
defparam \wb_csr_data[18] .is_wysiwyg = "true";
defparam \wb_csr_data[18] .power_up = "low";

cyclone10lp_lcell_comb \npc[18]~32 (
	.dataa(\pc_cntr[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[17]~31 ),
	.combout(\npc[18]~32_combout ),
	.cout(\npc[18]~33 ));
defparam \npc[18]~32 .lut_mask = 16'hA50A;
defparam \npc[18]~32 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~16 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[18]~32_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~16_combout ),
	.cout());
defparam \id_npc~16 .lut_mask = 16'h8080;
defparam \id_npc~16 .sum_lutc_input = "datac";

dffeas \id_npc[18] (
	.clk(clk_clk),
	.d(\id_npc~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[18]~q ),
	.prn(vcc));
defparam \id_npc[18] .is_wysiwyg = "true";
defparam \id_npc[18] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~16 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[18]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~16_combout ),
	.cout());
defparam \ex_npc~16 .lut_mask = 16'h8080;
defparam \ex_npc~16 .sum_lutc_input = "datac";

dffeas \ex_npc[18] (
	.clk(clk_clk),
	.d(\ex_npc~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[18]~q ),
	.prn(vcc));
defparam \ex_npc[18] .is_wysiwyg = "true";
defparam \ex_npc[18] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~14 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~14_combout ),
	.cout());
defparam \mem_npc~14 .lut_mask = 16'h8888;
defparam \mem_npc~14 .sum_lutc_input = "datac";

dffeas \mem_npc[18] (
	.clk(clk_clk),
	.d(\mem_npc~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[18]~q ),
	.prn(vcc));
defparam \mem_npc[18] .is_wysiwyg = "true";
defparam \mem_npc[18] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~14 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~14_combout ),
	.cout());
defparam \wb_npc~14 .lut_mask = 16'h8888;
defparam \wb_npc~14 .sum_lutc_input = "datac";

dffeas \wb_npc[18] (
	.clk(clk_clk),
	.d(\wb_npc~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[18]~q ),
	.prn(vcc));
defparam \wb_npc[18] .is_wysiwyg = "true";
defparam \wb_npc[18] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~16 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~16_combout ),
	.cout());
defparam \wb_alu_out~16 .lut_mask = 16'h8888;
defparam \wb_alu_out~16 .sum_lutc_input = "datac";

dffeas \wb_alu_out[18] (
	.clk(clk_clk),
	.d(\wb_alu_out~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[18]~q ),
	.prn(vcc));
defparam \wb_alu_out[18] .is_wysiwyg = "true";
defparam \wb_alu_out[18] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[18]~35 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[18]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[18]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[18]~35_combout ),
	.cout());
defparam \_T_3543__T_3854_data[18]~35 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[18]~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~77 (
	.dataa(\wb_dmem_read_data~36_combout ),
	.datab(av_readdata_pre_18),
	.datac(\wb_dmem_read_data~23_combout ),
	.datad(\wb_dmem_read_data[22]~32_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~77_combout ),
	.cout());
defparam \wb_dmem_read_data~77 .lut_mask = 16'h00AE;
defparam \wb_dmem_read_data~77 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[18] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~77_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[18]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[18] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[18] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[18]~36 (
	.dataa(\wb_csr_data[18]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[18]~35_combout ),
	.datad(\wb_dmem_read_data[18]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[18]~36_combout ),
	.cout());
defparam \_T_3543__T_3854_data[18]~36 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[18]~36 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a14 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[18]~36_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_a_first_bit_number = 14;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_b_first_bit_number = 14;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a14 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~18 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a14~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~18_combout ),
	.cout());
defparam \ex_rs_1~18 .lut_mask = 16'h8888;
defparam \ex_rs_1~18 .sum_lutc_input = "datac";

dffeas \ex_rs_1[18] (
	.clk(clk_clk),
	.d(\ex_rs_1~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[18]~q ),
	.prn(vcc));
defparam \ex_rs_1[18] .is_wysiwyg = "true";
defparam \ex_rs_1[18] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[18]~67 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_18),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[18]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[18]~67_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[18]~67 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[18]~67 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[18]~68 (
	.dataa(\ex_rs_1[18]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[18]~67_combout ),
	.datad(\wb_csr_data[18]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[18]~68_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[18]~68 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[18]~68 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[18]~69 (
	.dataa(\mem_alu_out[18]~q ),
	.datab(\ex_reg_rs2_bypass[18]~68_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[18]~69_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[18]~69 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[18]~69 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[18]~70 (
	.dataa(\ex_reg_rs2_bypass[18]~69_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[18]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[18]~70_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[18]~70 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[18]~70 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[18]~82 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\alu_io_op2[18]~58_combout ),
	.datad(\ex_reg_rs2_bypass[18]~70_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[18]~82_combout ),
	.cout());
defparam \alu_io_op2[18]~82 .lut_mask = 16'hF8F0;
defparam \alu_io_op2[18]~82 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a14 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[18]~36_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a14_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_a_first_bit_number = 14;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_b_first_bit_number = 14;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a14 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~18 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a14~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~18_combout ),
	.cout());
defparam \ex_rs_0~18 .lut_mask = 16'h0080;
defparam \ex_rs_0~18 .sum_lutc_input = "datac";

dffeas \ex_rs_0[18] (
	.clk(clk_clk),
	.d(\ex_rs_0~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[18]~q ),
	.prn(vcc));
defparam \ex_rs_0[18] .is_wysiwyg = "true";
defparam \ex_rs_0[18] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[18]~74 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(av_readdata_pre_18),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\wb_alu_out[18]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[18]~74_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[18]~74 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[18]~74 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[18]~75 (
	.dataa(\ex_rs_0[18]~q ),
	.datab(\ex_reg_rs1_bypass[2]~138_combout ),
	.datac(\ex_reg_rs1_bypass[18]~74_combout ),
	.datad(\wb_csr_data[18]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[18]~75_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[18]~75 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[18]~75 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[18]~76 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[18]~75_combout ),
	.datad(\mem_csr_data[18]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[18]~76_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[18]~76 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[18]~76 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[18]~77 (
	.dataa(\ex_reg_rs1_bypass[18]~76_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[18]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[18]~77_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[18]~77 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[18]~77 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[18]~104 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[18]~q ),
	.datad(\ex_reg_rs1_bypass[18]~77_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[18]~104_combout ),
	.cout());
defparam \alu_io_op1[18]~104 .lut_mask = 16'h6240;
defparam \alu_io_op1[18]~104 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~75 (
	.dataa(\mem_alu_out[26]~2_combout ),
	.datab(\alu|_T_139[18]~combout ),
	.datac(\alu|LessThan0~0_combout ),
	.datad(\alu|ShiftRight0~209_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~75_combout ),
	.cout());
defparam \mem_alu_out~75 .lut_mask = 16'h5E0E;
defparam \mem_alu_out~75 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~76 (
	.dataa(\alu_io_op1[18]~104_combout ),
	.datab(\alu_io_op2[18]~82_combout ),
	.datac(\mem_alu_out~75_combout ),
	.datad(\mem_alu_out[26]~2_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~76_combout ),
	.cout());
defparam \mem_alu_out~76 .lut_mask = 16'h86F0;
defparam \mem_alu_out~76 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~77 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[18]~104_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~76_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~77_combout ),
	.cout());
defparam \mem_alu_out~77 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~77 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~78 (
	.dataa(\alu_io_op2[18]~82_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~77_combout ),
	.datad(\alu|ShiftRight0~249_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~78_combout ),
	.cout());
defparam \mem_alu_out~78 .lut_mask = 16'hF838;
defparam \mem_alu_out~78 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~79 (
	.dataa(\mem_alu_out~78_combout ),
	.datab(\alu|_T_3[18]~36_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~79_combout ),
	.cout());
defparam \mem_alu_out~79 .lut_mask = 16'h00AC;
defparam \mem_alu_out~79 .sum_lutc_input = "datac";

dffeas \mem_alu_out[18] (
	.clk(clk_clk),
	.d(\mem_alu_out~79_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[18]~q ),
	.prn(vcc));
defparam \mem_alu_out[18] .is_wysiwyg = "true";
defparam \mem_alu_out[18] .power_up = "low";

cyclone10lp_lcell_comb \pc_cntr~58 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(\mem_alu_out[18]~q ),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[18]~32_combout ),
	.cin(gnd),
	.combout(\pc_cntr~58_combout ),
	.cout());
defparam \pc_cntr~58 .lut_mask = 16'hDAD0;
defparam \pc_cntr~58 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~59 (
	.dataa(\_T_3862[18]~36_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~58_combout ),
	.datad(\csr|mepc[18]~q ),
	.cin(gnd),
	.combout(\pc_cntr~59_combout ),
	.cout());
defparam \pc_cntr~59 .lut_mask = 16'hF2C2;
defparam \pc_cntr~59 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~60 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~59_combout ),
	.datac(\csr|mtvec[18]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~60_combout ),
	.cout());
defparam \pc_cntr~60 .lut_mask = 16'h88A0;
defparam \pc_cntr~60 .sum_lutc_input = "datac";

dffeas \pc_cntr[18] (
	.clk(clk_clk),
	.d(\pc_cntr~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[18]~q ),
	.prn(vcc));
defparam \pc_cntr[18] .is_wysiwyg = "true";
defparam \pc_cntr[18] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~17 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[18]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~17_combout ),
	.cout());
defparam \id_pc~17 .lut_mask = 16'h8080;
defparam \id_pc~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~17 (
	.dataa(id_pc_19),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~17_combout ),
	.cout());
defparam \ex_pc~17 .lut_mask = 16'h8080;
defparam \ex_pc~17 .sum_lutc_input = "datac";

dffeas \ex_pc[19] (
	.clk(clk_clk),
	.d(\ex_pc~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[19]~q ),
	.prn(vcc));
defparam \ex_pc[19] .is_wysiwyg = "true";
defparam \ex_pc[19] .power_up = "low";

cyclone10lp_lcell_comb \npc[19]~34 (
	.dataa(\pc_cntr[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[18]~33 ),
	.combout(\npc[19]~34_combout ),
	.cout(\npc[19]~35 ));
defparam \npc[19]~34 .lut_mask = 16'h5A5F;
defparam \npc[19]~34 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~17 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[19]~34_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~17_combout ),
	.cout());
defparam \id_npc~17 .lut_mask = 16'h8080;
defparam \id_npc~17 .sum_lutc_input = "datac";

dffeas \id_npc[19] (
	.clk(clk_clk),
	.d(\id_npc~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[19]~q ),
	.prn(vcc));
defparam \id_npc[19] .is_wysiwyg = "true";
defparam \id_npc[19] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~17 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[19]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~17_combout ),
	.cout());
defparam \ex_npc~17 .lut_mask = 16'h8080;
defparam \ex_npc~17 .sum_lutc_input = "datac";

dffeas \ex_npc[19] (
	.clk(clk_clk),
	.d(\ex_npc~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[19]~q ),
	.prn(vcc));
defparam \ex_npc[19] .is_wysiwyg = "true";
defparam \ex_npc[19] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~15 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[19]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~15_combout ),
	.cout());
defparam \mem_npc~15 .lut_mask = 16'h8888;
defparam \mem_npc~15 .sum_lutc_input = "datac";

dffeas \mem_npc[19] (
	.clk(clk_clk),
	.d(\mem_npc~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[19]~q ),
	.prn(vcc));
defparam \mem_npc[19] .is_wysiwyg = "true";
defparam \mem_npc[19] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~15 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[19]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~15_combout ),
	.cout());
defparam \wb_npc~15 .lut_mask = 16'h8888;
defparam \wb_npc~15 .sum_lutc_input = "datac";

dffeas \wb_npc[19] (
	.clk(clk_clk),
	.d(\wb_npc~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[19]~q ),
	.prn(vcc));
defparam \wb_npc[19] .is_wysiwyg = "true";
defparam \wb_npc[19] .power_up = "low";

cyclone10lp_lcell_comb \mem_csr_data~24 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[19]~135_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~24_combout ),
	.cout());
defparam \mem_csr_data~24 .lut_mask = 16'h8888;
defparam \mem_csr_data~24 .sum_lutc_input = "datac";

dffeas \mem_csr_data[19] (
	.clk(clk_clk),
	.d(\mem_csr_data~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[19]~q ),
	.prn(vcc));
defparam \mem_csr_data[19] .is_wysiwyg = "true";
defparam \mem_csr_data[19] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~17 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[19]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~17_combout ),
	.cout());
defparam \wb_csr_data~17 .lut_mask = 16'h8888;
defparam \wb_csr_data~17 .sum_lutc_input = "datac";

dffeas \wb_csr_data[19] (
	.clk(clk_clk),
	.d(\wb_csr_data~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[19]~q ),
	.prn(vcc));
defparam \wb_csr_data[19] .is_wysiwyg = "true";
defparam \wb_csr_data[19] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~17 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[19]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~17_combout ),
	.cout());
defparam \wb_alu_out~17 .lut_mask = 16'h8888;
defparam \wb_alu_out~17 .sum_lutc_input = "datac";

dffeas \wb_alu_out[19] (
	.clk(clk_clk),
	.d(\wb_alu_out~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[19]~q ),
	.prn(vcc));
defparam \wb_alu_out[19] .is_wysiwyg = "true";
defparam \wb_alu_out[19] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[19]~37 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[19]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[19]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[19]~37_combout ),
	.cout());
defparam \_T_3543__T_3854_data[19]~37 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[19]~37 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~78 (
	.dataa(\wb_dmem_read_data~30_combout ),
	.datab(av_readdata_pre_19),
	.datac(\wb_dmem_read_data~23_combout ),
	.datad(\wb_dmem_read_data[22]~32_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~78_combout ),
	.cout());
defparam \wb_dmem_read_data~78 .lut_mask = 16'h00AE;
defparam \wb_dmem_read_data~78 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[19] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[19]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[19] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[19] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[19]~38 (
	.dataa(\wb_npc[19]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[19]~37_combout ),
	.datad(\wb_dmem_read_data[19]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[19]~38_combout ),
	.cout());
defparam \_T_3543__T_3854_data[19]~38 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[19]~38 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a13 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[19]~38_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a13_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_a_first_bit_number = 13;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_b_first_bit_number = 13;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a13 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~19 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a13~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~19_combout ),
	.cout());
defparam \ex_rs_0~19 .lut_mask = 16'h0080;
defparam \ex_rs_0~19 .sum_lutc_input = "datac";

dffeas \ex_rs_0[19] (
	.clk(clk_clk),
	.d(\ex_rs_0~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[19]~q ),
	.prn(vcc));
defparam \ex_rs_0[19] .is_wysiwyg = "true";
defparam \ex_rs_0[19] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[19]~78 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(\ex_rs_0[19]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\wb_alu_out[19]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[19]~78_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[19]~78 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[19]~78 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[19]~79 (
	.dataa(av_readdata_pre_19),
	.datab(\ex_reg_rs1_bypass[2]~7_combout ),
	.datac(\ex_reg_rs1_bypass[19]~78_combout ),
	.datad(\wb_csr_data[19]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[19]~79_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[19]~79 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[19]~79 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[19]~80 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[19]~79_combout ),
	.datad(\mem_csr_data[19]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[19]~80_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[19]~80 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[19]~80 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[19]~81 (
	.dataa(\ex_reg_rs1_bypass[19]~80_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[19]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[19]~81_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[19]~81 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[19]~81 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[19]~105 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[19]~q ),
	.datad(\ex_reg_rs1_bypass[19]~81_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[19]~105_combout ),
	.cout());
defparam \alu_io_op1[19]~105 .lut_mask = 16'h6240;
defparam \alu_io_op1[19]~105 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[19]~59 (
	.dataa(\ex_inst[19]~q ),
	.datab(\mem_imm~7_combout ),
	.datac(\_T_3579~combout ),
	.datad(\ex_ctrl_alu_op2.10~q ),
	.cin(gnd),
	.combout(\alu_io_op2[19]~59_combout ),
	.cout());
defparam \alu_io_op2[19]~59 .lut_mask = 16'h00AC;
defparam \alu_io_op2[19]~59 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a13 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[19]~38_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_a_first_bit_number = 13;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_b_first_bit_number = 13;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a13 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~19 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a13~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~19_combout ),
	.cout());
defparam \ex_rs_1~19 .lut_mask = 16'h8888;
defparam \ex_rs_1~19 .sum_lutc_input = "datac";

dffeas \ex_rs_1[19] (
	.clk(clk_clk),
	.d(\ex_rs_1~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[19]~q ),
	.prn(vcc));
defparam \ex_rs_1[19] .is_wysiwyg = "true";
defparam \ex_rs_1[19] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[19]~71 (
	.dataa(\ex_reg_rs2_bypass[7]~5_combout ),
	.datab(\ex_rs_1[19]~q ),
	.datac(\ex_reg_rs2_bypass[7]~4_combout ),
	.datad(\wb_alu_out[19]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[19]~71_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[19]~71 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[19]~71 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[19]~72 (
	.dataa(av_readdata_pre_19),
	.datab(\ex_reg_rs2_bypass[7]~5_combout ),
	.datac(\ex_reg_rs2_bypass[19]~71_combout ),
	.datad(\wb_csr_data[19]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[19]~72_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[19]~72 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[19]~72 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[19]~73 (
	.dataa(\mem_alu_out[19]~q ),
	.datab(\ex_reg_rs2_bypass[19]~72_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[19]~73_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[19]~73 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[19]~73 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[19]~74 (
	.dataa(\ex_reg_rs2_bypass[19]~73_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[19]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[19]~74_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[19]~74 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[19]~74 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[19]~93 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\alu_io_op2[19]~59_combout ),
	.datad(\ex_reg_rs2_bypass[19]~74_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[19]~93_combout ),
	.cout());
defparam \alu_io_op2[19]~93 .lut_mask = 16'hF8F0;
defparam \alu_io_op2[19]~93 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~80 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\alu|_T_123[19]~combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~203_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~80_combout ),
	.cout());
defparam \mem_alu_out~80 .lut_mask = 16'hDAD0;
defparam \mem_alu_out~80 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~81 (
	.dataa(\alu_io_op1[19]~105_combout ),
	.datab(\alu_io_op2[19]~93_combout ),
	.datac(\mem_alu_out~80_combout ),
	.datad(\alu|LessThan0~0_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~81_combout ),
	.cout());
defparam \mem_alu_out~81 .lut_mask = 16'hF08E;
defparam \mem_alu_out~81 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~82 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[19]~93_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~81_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~82_combout ),
	.cout());
defparam \mem_alu_out~82 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~82 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~83 (
	.dataa(\alu_io_op1[19]~105_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~82_combout ),
	.datad(\alu|ShiftRight0~198_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~83_combout ),
	.cout());
defparam \mem_alu_out~83 .lut_mask = 16'hF838;
defparam \mem_alu_out~83 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~84 (
	.dataa(\mem_alu_out~83_combout ),
	.datab(\alu|_T_3[19]~38_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~84_combout ),
	.cout());
defparam \mem_alu_out~84 .lut_mask = 16'h00AC;
defparam \mem_alu_out~84 .sum_lutc_input = "datac";

dffeas \mem_alu_out[19] (
	.clk(clk_clk),
	.d(\mem_alu_out~84_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[19]~q ),
	.prn(vcc));
defparam \mem_alu_out[19] .is_wysiwyg = "true";
defparam \mem_alu_out[19] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~17 (
	.dataa(\ex_pc[19]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~17_combout ),
	.cout());
defparam \mem_pc~17 .lut_mask = 16'h8888;
defparam \mem_pc~17 .sum_lutc_input = "datac";

dffeas \mem_pc[19] (
	.clk(clk_clk),
	.d(\mem_pc~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[19]~q ),
	.prn(vcc));
defparam \mem_pc[19] .is_wysiwyg = "true";
defparam \mem_pc[19] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~34 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_inst[19]~q ),
	.datac(\mem_imm~7_combout ),
	.datad(\_T_3579~combout ),
	.cin(gnd),
	.combout(\mem_imm~34_combout ),
	.cout());
defparam \mem_imm~34 .lut_mask = 16'h88A0;
defparam \mem_imm~34 .sum_lutc_input = "datac";

dffeas \mem_imm[19] (
	.clk(clk_clk),
	.d(\mem_imm~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[19]~q ),
	.prn(vcc));
defparam \mem_imm[19] .is_wysiwyg = "true";
defparam \mem_imm[19] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[19]~38 (
	.dataa(\mem_pc[19]~q ),
	.datab(\mem_imm[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[18]~37 ),
	.combout(\_T_3862[19]~38_combout ),
	.cout(\_T_3862[19]~39 ));
defparam \_T_3862[19]~38 .lut_mask = 16'h9617;
defparam \_T_3862[19]~38 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~61 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[19]~38_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[19]~34_combout ),
	.cin(gnd),
	.combout(\pc_cntr~61_combout ),
	.cout());
defparam \pc_cntr~61 .lut_mask = 16'h5E0E;
defparam \pc_cntr~61 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~62 (
	.dataa(\mem_alu_out[19]~q ),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~61_combout ),
	.datad(\csr|mepc[19]~q ),
	.cin(gnd),
	.combout(\pc_cntr~62_combout ),
	.cout());
defparam \pc_cntr~62 .lut_mask = 16'hF838;
defparam \pc_cntr~62 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~63 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~62_combout ),
	.datac(\csr|mtvec[19]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~63_combout ),
	.cout());
defparam \pc_cntr~63 .lut_mask = 16'h88A0;
defparam \pc_cntr~63 .sum_lutc_input = "datac";

dffeas \pc_cntr[19] (
	.clk(clk_clk),
	.d(\pc_cntr~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[19]~q ),
	.prn(vcc));
defparam \pc_cntr[19] .is_wysiwyg = "true";
defparam \pc_cntr[19] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~18 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[19]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~18_combout ),
	.cout());
defparam \id_pc~18 .lut_mask = 16'h8080;
defparam \id_pc~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~18 (
	.dataa(id_pc_20),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~18_combout ),
	.cout());
defparam \ex_pc~18 .lut_mask = 16'h8080;
defparam \ex_pc~18 .sum_lutc_input = "datac";

dffeas \ex_pc[20] (
	.clk(clk_clk),
	.d(\ex_pc~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[20]~q ),
	.prn(vcc));
defparam \ex_pc[20] .is_wysiwyg = "true";
defparam \ex_pc[20] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~18 (
	.dataa(\ex_pc[20]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~18_combout ),
	.cout());
defparam \mem_pc~18 .lut_mask = 16'h8888;
defparam \mem_pc~18 .sum_lutc_input = "datac";

dffeas \mem_pc[20] (
	.clk(clk_clk),
	.d(\mem_pc~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[20]~q ),
	.prn(vcc));
defparam \mem_pc[20] .is_wysiwyg = "true";
defparam \mem_pc[20] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~9 (
	.dataa(\ex_csr_addr[0]~q ),
	.datab(\ex_ctrl_imm_type.011~q ),
	.datac(\ex_csr_addr[11]~q ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\mem_imm~9_combout ),
	.cout());
defparam \mem_imm~9 .lut_mask = 16'h88B8;
defparam \mem_imm~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~35 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\mem_imm~9_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_imm~35_combout ),
	.cout());
defparam \mem_imm~35 .lut_mask = 16'h8888;
defparam \mem_imm~35 .sum_lutc_input = "datac";

dffeas \mem_imm[20] (
	.clk(clk_clk),
	.d(\mem_imm~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[20]~q ),
	.prn(vcc));
defparam \mem_imm[20] .is_wysiwyg = "true";
defparam \mem_imm[20] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[20]~40 (
	.dataa(\mem_pc[20]~q ),
	.datab(\mem_imm[20]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[19]~39 ),
	.combout(\_T_3862[20]~40_combout ),
	.cout(\_T_3862[20]~41 ));
defparam \_T_3862[20]~40 .lut_mask = 16'h698E;
defparam \_T_3862[20]~40 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \mem_csr_data~31 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[20]~188_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~31_combout ),
	.cout());
defparam \mem_csr_data~31 .lut_mask = 16'h8888;
defparam \mem_csr_data~31 .sum_lutc_input = "datac";

dffeas \mem_csr_data[20] (
	.clk(clk_clk),
	.d(\mem_csr_data~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[20]~q ),
	.prn(vcc));
defparam \mem_csr_data[20] .is_wysiwyg = "true";
defparam \mem_csr_data[20] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~24 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~24_combout ),
	.cout());
defparam \wb_csr_data~24 .lut_mask = 16'h8888;
defparam \wb_csr_data~24 .sum_lutc_input = "datac";

dffeas \wb_csr_data[20] (
	.clk(clk_clk),
	.d(\wb_csr_data~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[20]~q ),
	.prn(vcc));
defparam \wb_csr_data[20] .is_wysiwyg = "true";
defparam \wb_csr_data[20] .power_up = "low";

cyclone10lp_lcell_comb \npc[20]~36 (
	.dataa(\pc_cntr[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[19]~35 ),
	.combout(\npc[20]~36_combout ),
	.cout(\npc[20]~37 ));
defparam \npc[20]~36 .lut_mask = 16'hA50A;
defparam \npc[20]~36 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~24 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[20]~36_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~24_combout ),
	.cout());
defparam \id_npc~24 .lut_mask = 16'h8080;
defparam \id_npc~24 .sum_lutc_input = "datac";

dffeas \id_npc[20] (
	.clk(clk_clk),
	.d(\id_npc~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[20]~q ),
	.prn(vcc));
defparam \id_npc[20] .is_wysiwyg = "true";
defparam \id_npc[20] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~24 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[20]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~24_combout ),
	.cout());
defparam \ex_npc~24 .lut_mask = 16'h8080;
defparam \ex_npc~24 .sum_lutc_input = "datac";

dffeas \ex_npc[20] (
	.clk(clk_clk),
	.d(\ex_npc~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[20]~q ),
	.prn(vcc));
defparam \ex_npc[20] .is_wysiwyg = "true";
defparam \ex_npc[20] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~22 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~22_combout ),
	.cout());
defparam \mem_npc~22 .lut_mask = 16'h8888;
defparam \mem_npc~22 .sum_lutc_input = "datac";

dffeas \mem_npc[20] (
	.clk(clk_clk),
	.d(\mem_npc~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[20]~q ),
	.prn(vcc));
defparam \mem_npc[20] .is_wysiwyg = "true";
defparam \mem_npc[20] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~22 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~22_combout ),
	.cout());
defparam \wb_npc~22 .lut_mask = 16'h8888;
defparam \wb_npc~22 .sum_lutc_input = "datac";

dffeas \wb_npc[20] (
	.clk(clk_clk),
	.d(\wb_npc~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[20]~q ),
	.prn(vcc));
defparam \wb_npc[20] .is_wysiwyg = "true";
defparam \wb_npc[20] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~24 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~24_combout ),
	.cout());
defparam \wb_alu_out~24 .lut_mask = 16'h8888;
defparam \wb_alu_out~24 .sum_lutc_input = "datac";

dffeas \wb_alu_out[20] (
	.clk(clk_clk),
	.d(\wb_alu_out~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[20]~q ),
	.prn(vcc));
defparam \wb_alu_out[20] .is_wysiwyg = "true";
defparam \wb_alu_out[20] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[20]~51 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[20]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[20]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[20]~51_combout ),
	.cout());
defparam \_T_3543__T_3854_data[20]~51 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[20]~51 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~79 (
	.dataa(\wb_dmem_read_data~36_combout ),
	.datab(av_readdata_pre_20),
	.datac(\wb_dmem_read_data~23_combout ),
	.datad(\wb_dmem_read_data[22]~32_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~79_combout ),
	.cout());
defparam \wb_dmem_read_data~79 .lut_mask = 16'h00AE;
defparam \wb_dmem_read_data~79 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[20] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~79_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[20]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[20] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[20] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[20]~52 (
	.dataa(\wb_csr_data[20]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[20]~51_combout ),
	.datad(\wb_dmem_read_data[20]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[20]~52_combout ),
	.cout());
defparam \_T_3543__T_3854_data[20]~52 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[20]~52 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a12 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[20]~52_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_a_first_bit_number = 12;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_b_first_bit_number = 12;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a12 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~27 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a12~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~27_combout ),
	.cout());
defparam \ex_rs_1~27 .lut_mask = 16'h8888;
defparam \ex_rs_1~27 .sum_lutc_input = "datac";

dffeas \ex_rs_1[20] (
	.clk(clk_clk),
	.d(\ex_rs_1~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[20]~q ),
	.prn(vcc));
defparam \ex_rs_1[20] .is_wysiwyg = "true";
defparam \ex_rs_1[20] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[20]~96 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_20),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[20]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[20]~96_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[20]~96 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[20]~96 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[20]~97 (
	.dataa(\ex_rs_1[20]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[20]~96_combout ),
	.datad(\wb_csr_data[20]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[20]~97_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[20]~97 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[20]~97 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[20]~98 (
	.dataa(\mem_alu_out[20]~q ),
	.datab(\ex_reg_rs2_bypass[20]~97_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[20]~98_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[20]~98 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[20]~98 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[20]~99 (
	.dataa(\ex_reg_rs2_bypass[20]~98_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[20]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[20]~99_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[20]~99 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[20]~99 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[20]~84 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_reg_rs2_bypass[20]~99_combout ),
	.datad(\mem_imm~9_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[20]~84_combout ),
	.cout());
defparam \alu_io_op2[20]~84 .lut_mask = 16'hB380;
defparam \alu_io_op2[20]~84 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a12 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[20]~52_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a12_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_a_first_bit_number = 12;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_b_first_bit_number = 12;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a12 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~26 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a12~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~26_combout ),
	.cout());
defparam \ex_rs_0~26 .lut_mask = 16'h0080;
defparam \ex_rs_0~26 .sum_lutc_input = "datac";

dffeas \ex_rs_0[20] (
	.clk(clk_clk),
	.d(\ex_rs_0~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[20]~q ),
	.prn(vcc));
defparam \ex_rs_0[20] .is_wysiwyg = "true";
defparam \ex_rs_0[20] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[20]~106 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(av_readdata_pre_20),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\wb_alu_out[20]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[20]~106_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[20]~106 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[20]~106 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[20]~107 (
	.dataa(\ex_rs_0[20]~q ),
	.datab(\ex_reg_rs1_bypass[2]~138_combout ),
	.datac(\ex_reg_rs1_bypass[20]~106_combout ),
	.datad(\wb_csr_data[20]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[20]~107_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[20]~107 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[20]~107 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[20]~108 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[20]~107_combout ),
	.datad(\mem_csr_data[20]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[20]~108_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[20]~108 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[20]~108 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[20]~109 (
	.dataa(\ex_reg_rs1_bypass[20]~108_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[20]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[20]~109_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[20]~109 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[20]~109 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[20]~112 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[20]~q ),
	.datad(\ex_reg_rs1_bypass[20]~109_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[20]~112_combout ),
	.cout());
defparam \alu_io_op1[20]~112 .lut_mask = 16'h6240;
defparam \alu_io_op1[20]~112 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~137 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\alu_io_op2[20]~84_combout ),
	.datad(\alu_io_op1[20]~112_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~137_combout ),
	.cout());
defparam \mem_alu_out~137 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~137 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~138 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~137_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~197_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~138_combout ),
	.cout());
defparam \mem_alu_out~138 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~138 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~99 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[20]~112_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~138_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~99_combout ),
	.cout());
defparam \mem_alu_out~99 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~99 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~100 (
	.dataa(\alu_io_op2[20]~84_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~99_combout ),
	.datad(\alu|ShiftRight0~195_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~100_combout ),
	.cout());
defparam \mem_alu_out~100 .lut_mask = 16'hF838;
defparam \mem_alu_out~100 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~101 (
	.dataa(\mem_alu_out~100_combout ),
	.datab(\alu|_T_3[20]~40_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~101_combout ),
	.cout());
defparam \mem_alu_out~101 .lut_mask = 16'h00AC;
defparam \mem_alu_out~101 .sum_lutc_input = "datac";

dffeas \mem_alu_out[20] (
	.clk(clk_clk),
	.d(\mem_alu_out~101_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[20]~q ),
	.prn(vcc));
defparam \mem_alu_out[20] .is_wysiwyg = "true";
defparam \mem_alu_out[20] .power_up = "low";

cyclone10lp_lcell_comb \pc_cntr~64 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(\mem_alu_out[20]~q ),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[20]~36_combout ),
	.cin(gnd),
	.combout(\pc_cntr~64_combout ),
	.cout());
defparam \pc_cntr~64 .lut_mask = 16'hDAD0;
defparam \pc_cntr~64 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~65 (
	.dataa(\_T_3862[20]~40_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~64_combout ),
	.datad(\csr|mepc[20]~q ),
	.cin(gnd),
	.combout(\pc_cntr~65_combout ),
	.cout());
defparam \pc_cntr~65 .lut_mask = 16'hF2C2;
defparam \pc_cntr~65 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~66 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~65_combout ),
	.datac(\csr|mtvec[20]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~66_combout ),
	.cout());
defparam \pc_cntr~66 .lut_mask = 16'h88A0;
defparam \pc_cntr~66 .sum_lutc_input = "datac";

dffeas \pc_cntr[20] (
	.clk(clk_clk),
	.d(\pc_cntr~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[20]~q ),
	.prn(vcc));
defparam \pc_cntr[20] .is_wysiwyg = "true";
defparam \pc_cntr[20] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~19 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[20]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~19_combout ),
	.cout());
defparam \id_pc~19 .lut_mask = 16'h8080;
defparam \id_pc~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~19 (
	.dataa(id_pc_21),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~19_combout ),
	.cout());
defparam \ex_pc~19 .lut_mask = 16'h8080;
defparam \ex_pc~19 .sum_lutc_input = "datac";

dffeas \ex_pc[21] (
	.clk(clk_clk),
	.d(\ex_pc~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[21]~q ),
	.prn(vcc));
defparam \ex_pc[21] .is_wysiwyg = "true";
defparam \ex_pc[21] .power_up = "low";

cyclone10lp_lcell_comb \npc[21]~38 (
	.dataa(\pc_cntr[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[20]~37 ),
	.combout(\npc[21]~38_combout ),
	.cout(\npc[21]~39 ));
defparam \npc[21]~38 .lut_mask = 16'h5A5F;
defparam \npc[21]~38 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~25 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[21]~38_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~25_combout ),
	.cout());
defparam \id_npc~25 .lut_mask = 16'h8080;
defparam \id_npc~25 .sum_lutc_input = "datac";

dffeas \id_npc[21] (
	.clk(clk_clk),
	.d(\id_npc~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[21]~q ),
	.prn(vcc));
defparam \id_npc[21] .is_wysiwyg = "true";
defparam \id_npc[21] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~25 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[21]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~25_combout ),
	.cout());
defparam \ex_npc~25 .lut_mask = 16'h8080;
defparam \ex_npc~25 .sum_lutc_input = "datac";

dffeas \ex_npc[21] (
	.clk(clk_clk),
	.d(\ex_npc~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[21]~q ),
	.prn(vcc));
defparam \ex_npc[21] .is_wysiwyg = "true";
defparam \ex_npc[21] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~23 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[21]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~23_combout ),
	.cout());
defparam \mem_npc~23 .lut_mask = 16'h8888;
defparam \mem_npc~23 .sum_lutc_input = "datac";

dffeas \mem_npc[21] (
	.clk(clk_clk),
	.d(\mem_npc~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[21]~q ),
	.prn(vcc));
defparam \mem_npc[21] .is_wysiwyg = "true";
defparam \mem_npc[21] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~23 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[21]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~23_combout ),
	.cout());
defparam \wb_npc~23 .lut_mask = 16'h8888;
defparam \wb_npc~23 .sum_lutc_input = "datac";

dffeas \wb_npc[21] (
	.clk(clk_clk),
	.d(\wb_npc~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[21]~q ),
	.prn(vcc));
defparam \wb_npc[21] .is_wysiwyg = "true";
defparam \wb_npc[21] .power_up = "low";

cyclone10lp_lcell_comb \mem_csr_data~37 (
	.dataa(\csr|io_out[21]~193_combout ),
	.datab(\csr|io_out[21]~194_combout ),
	.datac(\mem_ctrl_mem_wr~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~37_combout ),
	.cout());
defparam \mem_csr_data~37 .lut_mask = 16'hE0E0;
defparam \mem_csr_data~37 .sum_lutc_input = "datac";

dffeas \mem_csr_data[21] (
	.clk(clk_clk),
	.d(\mem_csr_data~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[21]~q ),
	.prn(vcc));
defparam \mem_csr_data[21] .is_wysiwyg = "true";
defparam \mem_csr_data[21] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~25 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[21]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~25_combout ),
	.cout());
defparam \wb_csr_data~25 .lut_mask = 16'h8888;
defparam \wb_csr_data~25 .sum_lutc_input = "datac";

dffeas \wb_csr_data[21] (
	.clk(clk_clk),
	.d(\wb_csr_data~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[21]~q ),
	.prn(vcc));
defparam \wb_csr_data[21] .is_wysiwyg = "true";
defparam \wb_csr_data[21] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~25 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[21]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~25_combout ),
	.cout());
defparam \wb_alu_out~25 .lut_mask = 16'h8888;
defparam \wb_alu_out~25 .sum_lutc_input = "datac";

dffeas \wb_alu_out[21] (
	.clk(clk_clk),
	.d(\wb_alu_out~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[21]~q ),
	.prn(vcc));
defparam \wb_alu_out[21] .is_wysiwyg = "true";
defparam \wb_alu_out[21] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[21]~53 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[21]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[21]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[21]~53_combout ),
	.cout());
defparam \_T_3543__T_3854_data[21]~53 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[21]~53 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~80 (
	.dataa(\wb_dmem_read_data~30_combout ),
	.datab(av_readdata_pre_21),
	.datac(\wb_dmem_read_data~23_combout ),
	.datad(\wb_dmem_read_data[22]~32_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~80_combout ),
	.cout());
defparam \wb_dmem_read_data~80 .lut_mask = 16'h00AE;
defparam \wb_dmem_read_data~80 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[21] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~80_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[21]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[21] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[21] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[21]~54 (
	.dataa(\wb_npc[21]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[21]~53_combout ),
	.datad(\wb_dmem_read_data[21]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[21]~54_combout ),
	.cout());
defparam \_T_3543__T_3854_data[21]~54 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[21]~54 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a11 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[21]~54_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a11_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_a_first_bit_number = 11;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_b_first_bit_number = 11;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a11 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~27 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a11~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~27_combout ),
	.cout());
defparam \ex_rs_0~27 .lut_mask = 16'h0080;
defparam \ex_rs_0~27 .sum_lutc_input = "datac";

dffeas \ex_rs_0[21] (
	.clk(clk_clk),
	.d(\ex_rs_0~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[21]~q ),
	.prn(vcc));
defparam \ex_rs_0[21] .is_wysiwyg = "true";
defparam \ex_rs_0[21] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[21]~110 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(\ex_rs_0[21]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\wb_alu_out[21]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[21]~110_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[21]~110 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[21]~110 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[21]~111 (
	.dataa(av_readdata_pre_21),
	.datab(\ex_reg_rs1_bypass[2]~7_combout ),
	.datac(\ex_reg_rs1_bypass[21]~110_combout ),
	.datad(\wb_csr_data[21]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[21]~111_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[21]~111 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[21]~111 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[21]~112 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[21]~111_combout ),
	.datad(\mem_csr_data[21]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[21]~112_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[21]~112 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[21]~112 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[21]~113 (
	.dataa(\ex_reg_rs1_bypass[21]~112_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[21]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[21]~113_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[21]~113 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[21]~113 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[21]~113 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[21]~q ),
	.datad(\ex_reg_rs1_bypass[21]~113_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[21]~113_combout ),
	.cout());
defparam \alu_io_op1[21]~113 .lut_mask = 16'h6240;
defparam \alu_io_op1[21]~113 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a11 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[21]~54_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_a_first_bit_number = 11;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_b_first_bit_number = 11;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a11 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~26 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a11~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~26_combout ),
	.cout());
defparam \ex_rs_1~26 .lut_mask = 16'h8888;
defparam \ex_rs_1~26 .sum_lutc_input = "datac";

dffeas \ex_rs_1[21] (
	.clk(clk_clk),
	.d(\ex_rs_1~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[21]~q ),
	.prn(vcc));
defparam \ex_rs_1[21] .is_wysiwyg = "true";
defparam \ex_rs_1[21] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[21]~92 (
	.dataa(\ex_reg_rs2_bypass[7]~5_combout ),
	.datab(\ex_rs_1[21]~q ),
	.datac(\ex_reg_rs2_bypass[7]~4_combout ),
	.datad(\wb_alu_out[21]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[21]~92_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[21]~92 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[21]~92 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[21]~93 (
	.dataa(av_readdata_pre_21),
	.datab(\ex_reg_rs2_bypass[7]~5_combout ),
	.datac(\ex_reg_rs2_bypass[21]~92_combout ),
	.datad(\wb_csr_data[21]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[21]~93_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[21]~93 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[21]~93 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[21]~94 (
	.dataa(\mem_alu_out[21]~q ),
	.datab(\ex_reg_rs2_bypass[21]~93_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[21]~94_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[21]~94 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[21]~94 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[21]~95 (
	.dataa(\ex_reg_rs2_bypass[21]~94_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[21]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[21]~95_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[21]~95 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[21]~95 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~8 (
	.dataa(\ex_csr_addr[1]~q ),
	.datab(\ex_ctrl_imm_type.011~q ),
	.datac(\ex_csr_addr[11]~q ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\mem_imm~8_combout ),
	.cout());
defparam \mem_imm~8 .lut_mask = 16'h88B8;
defparam \mem_imm~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[21]~83 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_reg_rs2_bypass[21]~95_combout ),
	.datad(\mem_imm~8_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[21]~83_combout ),
	.cout());
defparam \alu_io_op2[21]~83 .lut_mask = 16'hB380;
defparam \alu_io_op2[21]~83 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~102 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\alu|_T_123[21]~combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~190_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~102_combout ),
	.cout());
defparam \mem_alu_out~102 .lut_mask = 16'hDAD0;
defparam \mem_alu_out~102 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~103 (
	.dataa(\alu_io_op1[21]~113_combout ),
	.datab(\alu_io_op2[21]~83_combout ),
	.datac(\mem_alu_out~102_combout ),
	.datad(\alu|LessThan0~0_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~103_combout ),
	.cout());
defparam \mem_alu_out~103 .lut_mask = 16'hF08E;
defparam \mem_alu_out~103 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~104 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[21]~83_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~103_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~104_combout ),
	.cout());
defparam \mem_alu_out~104 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~104 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~105 (
	.dataa(\alu_io_op1[21]~113_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~104_combout ),
	.datad(\alu|ShiftRight0~188_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~105_combout ),
	.cout());
defparam \mem_alu_out~105 .lut_mask = 16'hF838;
defparam \mem_alu_out~105 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~106 (
	.dataa(\mem_alu_out~105_combout ),
	.datab(\alu|_T_3[21]~42_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~106_combout ),
	.cout());
defparam \mem_alu_out~106 .lut_mask = 16'h00AC;
defparam \mem_alu_out~106 .sum_lutc_input = "datac";

dffeas \mem_alu_out[21] (
	.clk(clk_clk),
	.d(\mem_alu_out~106_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[21]~q ),
	.prn(vcc));
defparam \mem_alu_out[21] .is_wysiwyg = "true";
defparam \mem_alu_out[21] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~19 (
	.dataa(\ex_pc[21]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~19_combout ),
	.cout());
defparam \mem_pc~19 .lut_mask = 16'h8888;
defparam \mem_pc~19 .sum_lutc_input = "datac";

dffeas \mem_pc[21] (
	.clk(clk_clk),
	.d(\mem_pc~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[21]~q ),
	.prn(vcc));
defparam \mem_pc[21] .is_wysiwyg = "true";
defparam \mem_pc[21] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~36 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\mem_imm~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_imm~36_combout ),
	.cout());
defparam \mem_imm~36 .lut_mask = 16'h8888;
defparam \mem_imm~36 .sum_lutc_input = "datac";

dffeas \mem_imm[21] (
	.clk(clk_clk),
	.d(\mem_imm~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[21]~q ),
	.prn(vcc));
defparam \mem_imm[21] .is_wysiwyg = "true";
defparam \mem_imm[21] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[21]~42 (
	.dataa(\mem_pc[21]~q ),
	.datab(\mem_imm[21]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[20]~41 ),
	.combout(\_T_3862[21]~42_combout ),
	.cout(\_T_3862[21]~43 ));
defparam \_T_3862[21]~42 .lut_mask = 16'h9617;
defparam \_T_3862[21]~42 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~67 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[21]~42_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[21]~38_combout ),
	.cin(gnd),
	.combout(\pc_cntr~67_combout ),
	.cout());
defparam \pc_cntr~67 .lut_mask = 16'h5E0E;
defparam \pc_cntr~67 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~68 (
	.dataa(\mem_alu_out[21]~q ),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~67_combout ),
	.datad(\csr|mepc[21]~q ),
	.cin(gnd),
	.combout(\pc_cntr~68_combout ),
	.cout());
defparam \pc_cntr~68 .lut_mask = 16'hF838;
defparam \pc_cntr~68 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~69 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~68_combout ),
	.datac(\csr|mtvec[21]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~69_combout ),
	.cout());
defparam \pc_cntr~69 .lut_mask = 16'h88A0;
defparam \pc_cntr~69 .sum_lutc_input = "datac";

dffeas \pc_cntr[21] (
	.clk(clk_clk),
	.d(\pc_cntr~69_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[21]~q ),
	.prn(vcc));
defparam \pc_cntr[21] .is_wysiwyg = "true";
defparam \pc_cntr[21] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~20 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[21]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~20_combout ),
	.cout());
defparam \id_pc~20 .lut_mask = 16'h8080;
defparam \id_pc~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~20 (
	.dataa(id_pc_22),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~20_combout ),
	.cout());
defparam \ex_pc~20 .lut_mask = 16'h8080;
defparam \ex_pc~20 .sum_lutc_input = "datac";

dffeas \ex_pc[22] (
	.clk(clk_clk),
	.d(\ex_pc~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[22]~q ),
	.prn(vcc));
defparam \ex_pc[22] .is_wysiwyg = "true";
defparam \ex_pc[22] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~20 (
	.dataa(\ex_pc[22]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~20_combout ),
	.cout());
defparam \mem_pc~20 .lut_mask = 16'h8888;
defparam \mem_pc~20 .sum_lutc_input = "datac";

dffeas \mem_pc[22] (
	.clk(clk_clk),
	.d(\mem_pc~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[22]~q ),
	.prn(vcc));
defparam \mem_pc[22] .is_wysiwyg = "true";
defparam \mem_pc[22] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~10 (
	.dataa(\ex_csr_addr[2]~q ),
	.datab(\ex_ctrl_imm_type.011~q ),
	.datac(\ex_csr_addr[11]~q ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\mem_imm~10_combout ),
	.cout());
defparam \mem_imm~10 .lut_mask = 16'h88B8;
defparam \mem_imm~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~37 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\mem_imm~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_imm~37_combout ),
	.cout());
defparam \mem_imm~37 .lut_mask = 16'h8888;
defparam \mem_imm~37 .sum_lutc_input = "datac";

dffeas \mem_imm[22] (
	.clk(clk_clk),
	.d(\mem_imm~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[22]~q ),
	.prn(vcc));
defparam \mem_imm[22] .is_wysiwyg = "true";
defparam \mem_imm[22] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[22]~44 (
	.dataa(\mem_pc[22]~q ),
	.datab(\mem_imm[22]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[21]~43 ),
	.combout(\_T_3862[22]~44_combout ),
	.cout(\_T_3862[22]~45 ));
defparam \_T_3862[22]~44 .lut_mask = 16'h698E;
defparam \_T_3862[22]~44 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \mem_csr_data~32 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[22]~202_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~32_combout ),
	.cout());
defparam \mem_csr_data~32 .lut_mask = 16'h8888;
defparam \mem_csr_data~32 .sum_lutc_input = "datac";

dffeas \mem_csr_data[22] (
	.clk(clk_clk),
	.d(\mem_csr_data~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[22]~q ),
	.prn(vcc));
defparam \mem_csr_data[22] .is_wysiwyg = "true";
defparam \mem_csr_data[22] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~26 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[22]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~26_combout ),
	.cout());
defparam \wb_csr_data~26 .lut_mask = 16'h8888;
defparam \wb_csr_data~26 .sum_lutc_input = "datac";

dffeas \wb_csr_data[22] (
	.clk(clk_clk),
	.d(\wb_csr_data~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[22]~q ),
	.prn(vcc));
defparam \wb_csr_data[22] .is_wysiwyg = "true";
defparam \wb_csr_data[22] .power_up = "low";

cyclone10lp_lcell_comb \npc[22]~40 (
	.dataa(\pc_cntr[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[21]~39 ),
	.combout(\npc[22]~40_combout ),
	.cout(\npc[22]~41 ));
defparam \npc[22]~40 .lut_mask = 16'hA50A;
defparam \npc[22]~40 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~26 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[22]~40_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~26_combout ),
	.cout());
defparam \id_npc~26 .lut_mask = 16'h8080;
defparam \id_npc~26 .sum_lutc_input = "datac";

dffeas \id_npc[22] (
	.clk(clk_clk),
	.d(\id_npc~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[22]~q ),
	.prn(vcc));
defparam \id_npc[22] .is_wysiwyg = "true";
defparam \id_npc[22] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~26 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[22]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~26_combout ),
	.cout());
defparam \ex_npc~26 .lut_mask = 16'h8080;
defparam \ex_npc~26 .sum_lutc_input = "datac";

dffeas \ex_npc[22] (
	.clk(clk_clk),
	.d(\ex_npc~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[22]~q ),
	.prn(vcc));
defparam \ex_npc[22] .is_wysiwyg = "true";
defparam \ex_npc[22] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~24 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[22]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~24_combout ),
	.cout());
defparam \mem_npc~24 .lut_mask = 16'h8888;
defparam \mem_npc~24 .sum_lutc_input = "datac";

dffeas \mem_npc[22] (
	.clk(clk_clk),
	.d(\mem_npc~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[22]~q ),
	.prn(vcc));
defparam \mem_npc[22] .is_wysiwyg = "true";
defparam \mem_npc[22] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~24 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[22]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~24_combout ),
	.cout());
defparam \wb_npc~24 .lut_mask = 16'h8888;
defparam \wb_npc~24 .sum_lutc_input = "datac";

dffeas \wb_npc[22] (
	.clk(clk_clk),
	.d(\wb_npc~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[22]~q ),
	.prn(vcc));
defparam \wb_npc[22] .is_wysiwyg = "true";
defparam \wb_npc[22] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~26 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[22]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~26_combout ),
	.cout());
defparam \wb_alu_out~26 .lut_mask = 16'h8888;
defparam \wb_alu_out~26 .sum_lutc_input = "datac";

dffeas \wb_alu_out[22] (
	.clk(clk_clk),
	.d(\wb_alu_out~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[22]~q ),
	.prn(vcc));
defparam \wb_alu_out[22] .is_wysiwyg = "true";
defparam \wb_alu_out[22] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[22]~55 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[22]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[22]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[22]~55_combout ),
	.cout());
defparam \_T_3543__T_3854_data[22]~55 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[22]~55 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~81 (
	.dataa(\wb_dmem_read_data~36_combout ),
	.datab(av_readdata_pre_22),
	.datac(\wb_dmem_read_data~23_combout ),
	.datad(\wb_dmem_read_data[22]~32_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~81_combout ),
	.cout());
defparam \wb_dmem_read_data~81 .lut_mask = 16'h00AE;
defparam \wb_dmem_read_data~81 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[22] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~81_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[22]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[22] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[22] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[22]~56 (
	.dataa(\wb_csr_data[22]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[22]~55_combout ),
	.datad(\wb_dmem_read_data[22]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[22]~56_combout ),
	.cout());
defparam \_T_3543__T_3854_data[22]~56 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[22]~56 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a10 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[22]~56_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_a_first_bit_number = 10;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_b_first_bit_number = 10;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a10 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~28 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a10~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~28_combout ),
	.cout());
defparam \ex_rs_1~28 .lut_mask = 16'h8888;
defparam \ex_rs_1~28 .sum_lutc_input = "datac";

dffeas \ex_rs_1[22] (
	.clk(clk_clk),
	.d(\ex_rs_1~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[22]~q ),
	.prn(vcc));
defparam \ex_rs_1[22] .is_wysiwyg = "true";
defparam \ex_rs_1[22] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[22]~100 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_22),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[22]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[22]~100_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[22]~100 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[22]~100 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[22]~101 (
	.dataa(\ex_rs_1[22]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[22]~100_combout ),
	.datad(\wb_csr_data[22]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[22]~101_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[22]~101 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[22]~101 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[22]~102 (
	.dataa(\mem_alu_out[22]~q ),
	.datab(\ex_reg_rs2_bypass[22]~101_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[22]~102_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[22]~102 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[22]~102 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[22]~103 (
	.dataa(\ex_reg_rs2_bypass[22]~102_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[22]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[22]~103_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[22]~103 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[22]~103 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[22]~85 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_reg_rs2_bypass[22]~103_combout ),
	.datad(\mem_imm~10_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[22]~85_combout ),
	.cout());
defparam \alu_io_op2[22]~85 .lut_mask = 16'hB380;
defparam \alu_io_op2[22]~85 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a10 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[22]~56_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a10_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_a_first_bit_number = 10;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_b_first_bit_number = 10;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a10 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~28 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a10~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~28_combout ),
	.cout());
defparam \ex_rs_0~28 .lut_mask = 16'h0080;
defparam \ex_rs_0~28 .sum_lutc_input = "datac";

dffeas \ex_rs_0[22] (
	.clk(clk_clk),
	.d(\ex_rs_0~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[22]~q ),
	.prn(vcc));
defparam \ex_rs_0[22] .is_wysiwyg = "true";
defparam \ex_rs_0[22] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[22]~114 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(av_readdata_pre_22),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\wb_alu_out[22]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[22]~114_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[22]~114 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[22]~114 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[22]~115 (
	.dataa(\ex_rs_0[22]~q ),
	.datab(\ex_reg_rs1_bypass[2]~138_combout ),
	.datac(\ex_reg_rs1_bypass[22]~114_combout ),
	.datad(\wb_csr_data[22]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[22]~115_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[22]~115 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[22]~115 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[22]~116 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[22]~115_combout ),
	.datad(\mem_csr_data[22]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[22]~116_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[22]~116 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[22]~116 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[22]~117 (
	.dataa(\ex_reg_rs1_bypass[22]~116_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[22]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[22]~117_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[22]~117 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[22]~117 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[22]~114 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[22]~q ),
	.datad(\ex_reg_rs1_bypass[22]~117_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[22]~114_combout ),
	.cout());
defparam \alu_io_op1[22]~114 .lut_mask = 16'h6240;
defparam \alu_io_op1[22]~114 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~135 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\alu_io_op2[22]~85_combout ),
	.datad(\alu_io_op1[22]~114_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~135_combout ),
	.cout());
defparam \mem_alu_out~135 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~135 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~136 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~135_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~183_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~136_combout ),
	.cout());
defparam \mem_alu_out~136 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~136 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~107 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[22]~114_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~136_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~107_combout ),
	.cout());
defparam \mem_alu_out~107 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~107 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~108 (
	.dataa(\alu_io_op2[22]~85_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~107_combout ),
	.datad(\alu|ShiftRight0~180_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~108_combout ),
	.cout());
defparam \mem_alu_out~108 .lut_mask = 16'hF838;
defparam \mem_alu_out~108 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~109 (
	.dataa(\mem_alu_out~108_combout ),
	.datab(\alu|_T_3[22]~44_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~109_combout ),
	.cout());
defparam \mem_alu_out~109 .lut_mask = 16'h00AC;
defparam \mem_alu_out~109 .sum_lutc_input = "datac";

dffeas \mem_alu_out[22] (
	.clk(clk_clk),
	.d(\mem_alu_out~109_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[22]~q ),
	.prn(vcc));
defparam \mem_alu_out[22] .is_wysiwyg = "true";
defparam \mem_alu_out[22] .power_up = "low";

cyclone10lp_lcell_comb \pc_cntr~70 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(\mem_alu_out[22]~q ),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[22]~40_combout ),
	.cin(gnd),
	.combout(\pc_cntr~70_combout ),
	.cout());
defparam \pc_cntr~70 .lut_mask = 16'hDAD0;
defparam \pc_cntr~70 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~71 (
	.dataa(\_T_3862[22]~44_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~70_combout ),
	.datad(\csr|mepc[22]~q ),
	.cin(gnd),
	.combout(\pc_cntr~71_combout ),
	.cout());
defparam \pc_cntr~71 .lut_mask = 16'hF2C2;
defparam \pc_cntr~71 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~72 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~71_combout ),
	.datac(\csr|mtvec[22]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~72_combout ),
	.cout());
defparam \pc_cntr~72 .lut_mask = 16'h88A0;
defparam \pc_cntr~72 .sum_lutc_input = "datac";

dffeas \pc_cntr[22] (
	.clk(clk_clk),
	.d(\pc_cntr~72_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[22]~q ),
	.prn(vcc));
defparam \pc_cntr[22] .is_wysiwyg = "true";
defparam \pc_cntr[22] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~21 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[22]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~21_combout ),
	.cout());
defparam \id_pc~21 .lut_mask = 16'h8080;
defparam \id_pc~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~21 (
	.dataa(id_pc_23),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~21_combout ),
	.cout());
defparam \ex_pc~21 .lut_mask = 16'h8080;
defparam \ex_pc~21 .sum_lutc_input = "datac";

dffeas \ex_pc[23] (
	.clk(clk_clk),
	.d(\ex_pc~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[23]~q ),
	.prn(vcc));
defparam \ex_pc[23] .is_wysiwyg = "true";
defparam \ex_pc[23] .power_up = "low";

cyclone10lp_lcell_comb \npc[23]~42 (
	.dataa(\pc_cntr[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[22]~41 ),
	.combout(\npc[23]~42_combout ),
	.cout(\npc[23]~43 ));
defparam \npc[23]~42 .lut_mask = 16'h5A5F;
defparam \npc[23]~42 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~27 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[23]~42_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~27_combout ),
	.cout());
defparam \id_npc~27 .lut_mask = 16'h8080;
defparam \id_npc~27 .sum_lutc_input = "datac";

dffeas \id_npc[23] (
	.clk(clk_clk),
	.d(\id_npc~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[23]~q ),
	.prn(vcc));
defparam \id_npc[23] .is_wysiwyg = "true";
defparam \id_npc[23] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~27 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[23]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~27_combout ),
	.cout());
defparam \ex_npc~27 .lut_mask = 16'h8080;
defparam \ex_npc~27 .sum_lutc_input = "datac";

dffeas \ex_npc[23] (
	.clk(clk_clk),
	.d(\ex_npc~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[23]~q ),
	.prn(vcc));
defparam \ex_npc[23] .is_wysiwyg = "true";
defparam \ex_npc[23] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~25 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[23]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~25_combout ),
	.cout());
defparam \mem_npc~25 .lut_mask = 16'h8888;
defparam \mem_npc~25 .sum_lutc_input = "datac";

dffeas \mem_npc[23] (
	.clk(clk_clk),
	.d(\mem_npc~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[23]~q ),
	.prn(vcc));
defparam \mem_npc[23] .is_wysiwyg = "true";
defparam \mem_npc[23] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~25 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[23]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~25_combout ),
	.cout());
defparam \wb_npc~25 .lut_mask = 16'h8888;
defparam \wb_npc~25 .sum_lutc_input = "datac";

dffeas \wb_npc[23] (
	.clk(clk_clk),
	.d(\wb_npc~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[23]~q ),
	.prn(vcc));
defparam \wb_npc[23] .is_wysiwyg = "true";
defparam \wb_npc[23] .power_up = "low";

cyclone10lp_lcell_comb \mem_csr_data~33 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[23]~209_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~33_combout ),
	.cout());
defparam \mem_csr_data~33 .lut_mask = 16'h8888;
defparam \mem_csr_data~33 .sum_lutc_input = "datac";

dffeas \mem_csr_data[23] (
	.clk(clk_clk),
	.d(\mem_csr_data~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[23]~q ),
	.prn(vcc));
defparam \mem_csr_data[23] .is_wysiwyg = "true";
defparam \mem_csr_data[23] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~27 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[23]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~27_combout ),
	.cout());
defparam \wb_csr_data~27 .lut_mask = 16'h8888;
defparam \wb_csr_data~27 .sum_lutc_input = "datac";

dffeas \wb_csr_data[23] (
	.clk(clk_clk),
	.d(\wb_csr_data~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[23]~q ),
	.prn(vcc));
defparam \wb_csr_data[23] .is_wysiwyg = "true";
defparam \wb_csr_data[23] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~27 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[23]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~27_combout ),
	.cout());
defparam \wb_alu_out~27 .lut_mask = 16'h8888;
defparam \wb_alu_out~27 .sum_lutc_input = "datac";

dffeas \wb_alu_out[23] (
	.clk(clk_clk),
	.d(\wb_alu_out~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[23]~q ),
	.prn(vcc));
defparam \wb_alu_out[23] .is_wysiwyg = "true";
defparam \wb_alu_out[23] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[23]~57 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[23]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[23]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[23]~57_combout ),
	.cout());
defparam \_T_3543__T_3854_data[23]~57 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[23]~57 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~82 (
	.dataa(av_readdata_pre_31),
	.datab(av_readdata_pre_15),
	.datac(mem_alu_out_1),
	.datad(mem_alu_out_0),
	.cin(gnd),
	.combout(\wb_dmem_read_data~82_combout ),
	.cout());
defparam \wb_dmem_read_data~82 .lut_mask = 16'h00AC;
defparam \wb_dmem_read_data~82 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~83 (
	.dataa(mem_ctrl_mem_wr01),
	.datab(\wb_dmem_read_data~39_combout ),
	.datac(Equal73),
	.datad(\wb_dmem_read_data~82_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~83_combout ),
	.cout());
defparam \wb_dmem_read_data~83 .lut_mask = 16'hA888;
defparam \wb_dmem_read_data~83 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~84 (
	.dataa(\wb_dmem_read_data~83_combout ),
	.datab(av_readdata_pre_23),
	.datac(gnd),
	.datad(\wb_dmem_read_data~23_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~84_combout ),
	.cout());
defparam \wb_dmem_read_data~84 .lut_mask = 16'hAAEE;
defparam \wb_dmem_read_data~84 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[23] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~84_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[23]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[23] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[23] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[23]~58 (
	.dataa(\wb_npc[23]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[23]~57_combout ),
	.datad(\wb_dmem_read_data[23]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[23]~58_combout ),
	.cout());
defparam \_T_3543__T_3854_data[23]~58 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[23]~58 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a9 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[23]~58_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a9_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_a_first_bit_number = 9;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_b_first_bit_number = 9;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a9 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~29 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a9~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~29_combout ),
	.cout());
defparam \ex_rs_0~29 .lut_mask = 16'h0080;
defparam \ex_rs_0~29 .sum_lutc_input = "datac";

dffeas \ex_rs_0[23] (
	.clk(clk_clk),
	.d(\ex_rs_0~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[23]~q ),
	.prn(vcc));
defparam \ex_rs_0[23] .is_wysiwyg = "true";
defparam \ex_rs_0[23] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[23]~118 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(\ex_rs_0[23]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\wb_alu_out[23]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[23]~118_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[23]~118 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[23]~118 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[23]~119 (
	.dataa(av_readdata_pre_23),
	.datab(\ex_reg_rs1_bypass[2]~7_combout ),
	.datac(\ex_reg_rs1_bypass[23]~118_combout ),
	.datad(\wb_csr_data[23]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[23]~119_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[23]~119 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[23]~119 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[23]~120 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[23]~119_combout ),
	.datad(\mem_csr_data[23]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[23]~120_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[23]~120 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[23]~120 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[23]~121 (
	.dataa(\ex_reg_rs1_bypass[23]~120_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[23]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[23]~121_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[23]~121 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[23]~121 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[23]~119 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[23]~q ),
	.datad(\ex_reg_rs1_bypass[23]~121_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[23]~119_combout ),
	.cout());
defparam \alu_io_op1[23]~119 .lut_mask = 16'h6240;
defparam \alu_io_op1[23]~119 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a9 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[23]~58_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_a_first_bit_number = 9;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_b_first_bit_number = 9;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a9 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~29 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a9~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~29_combout ),
	.cout());
defparam \ex_rs_1~29 .lut_mask = 16'h8888;
defparam \ex_rs_1~29 .sum_lutc_input = "datac";

dffeas \ex_rs_1[23] (
	.clk(clk_clk),
	.d(\ex_rs_1~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[23]~q ),
	.prn(vcc));
defparam \ex_rs_1[23] .is_wysiwyg = "true";
defparam \ex_rs_1[23] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[23]~104 (
	.dataa(\ex_reg_rs2_bypass[7]~5_combout ),
	.datab(\ex_rs_1[23]~q ),
	.datac(\ex_reg_rs2_bypass[7]~4_combout ),
	.datad(\wb_alu_out[23]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[23]~104_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[23]~104 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[23]~104 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[23]~105 (
	.dataa(av_readdata_pre_23),
	.datab(\ex_reg_rs2_bypass[7]~5_combout ),
	.datac(\ex_reg_rs2_bypass[23]~104_combout ),
	.datad(\wb_csr_data[23]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[23]~105_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[23]~105 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[23]~105 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[23]~106 (
	.dataa(\mem_alu_out[23]~q ),
	.datab(\ex_reg_rs2_bypass[23]~105_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[23]~106_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[23]~106 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[23]~106 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[23]~107 (
	.dataa(\ex_reg_rs2_bypass[23]~106_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[23]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[23]~107_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[23]~107 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[23]~107 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~11 (
	.dataa(\ex_csr_addr[3]~q ),
	.datab(\ex_ctrl_imm_type.011~q ),
	.datac(\ex_csr_addr[11]~q ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\mem_imm~11_combout ),
	.cout());
defparam \mem_imm~11 .lut_mask = 16'h88B8;
defparam \mem_imm~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[23]~86 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_reg_rs2_bypass[23]~107_combout ),
	.datad(\mem_imm~11_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[23]~86_combout ),
	.cout());
defparam \alu_io_op2[23]~86 .lut_mask = 16'hB380;
defparam \alu_io_op2[23]~86 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~110 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\alu|_T_123[23]~combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~175_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~110_combout ),
	.cout());
defparam \mem_alu_out~110 .lut_mask = 16'hDAD0;
defparam \mem_alu_out~110 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~111 (
	.dataa(\alu_io_op1[23]~119_combout ),
	.datab(\alu_io_op2[23]~86_combout ),
	.datac(\mem_alu_out~110_combout ),
	.datad(\alu|LessThan0~0_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~111_combout ),
	.cout());
defparam \mem_alu_out~111 .lut_mask = 16'hF08E;
defparam \mem_alu_out~111 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~112 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[23]~86_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~111_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~112_combout ),
	.cout());
defparam \mem_alu_out~112 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~112 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~113 (
	.dataa(\alu_io_op1[23]~119_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~112_combout ),
	.datad(\alu|ShiftRight0~173_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~113_combout ),
	.cout());
defparam \mem_alu_out~113 .lut_mask = 16'hF838;
defparam \mem_alu_out~113 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~114 (
	.dataa(\mem_alu_out~113_combout ),
	.datab(\alu|_T_3[23]~46_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~114_combout ),
	.cout());
defparam \mem_alu_out~114 .lut_mask = 16'h00AC;
defparam \mem_alu_out~114 .sum_lutc_input = "datac";

dffeas \mem_alu_out[23] (
	.clk(clk_clk),
	.d(\mem_alu_out~114_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[23]~q ),
	.prn(vcc));
defparam \mem_alu_out[23] .is_wysiwyg = "true";
defparam \mem_alu_out[23] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~21 (
	.dataa(\ex_pc[23]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~21_combout ),
	.cout());
defparam \mem_pc~21 .lut_mask = 16'h8888;
defparam \mem_pc~21 .sum_lutc_input = "datac";

dffeas \mem_pc[23] (
	.clk(clk_clk),
	.d(\mem_pc~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[23]~q ),
	.prn(vcc));
defparam \mem_pc[23] .is_wysiwyg = "true";
defparam \mem_pc[23] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~38 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\mem_imm~11_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_imm~38_combout ),
	.cout());
defparam \mem_imm~38 .lut_mask = 16'h8888;
defparam \mem_imm~38 .sum_lutc_input = "datac";

dffeas \mem_imm[23] (
	.clk(clk_clk),
	.d(\mem_imm~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[23]~q ),
	.prn(vcc));
defparam \mem_imm[23] .is_wysiwyg = "true";
defparam \mem_imm[23] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[23]~46 (
	.dataa(\mem_pc[23]~q ),
	.datab(\mem_imm[23]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[22]~45 ),
	.combout(\_T_3862[23]~46_combout ),
	.cout(\_T_3862[23]~47 ));
defparam \_T_3862[23]~46 .lut_mask = 16'h9617;
defparam \_T_3862[23]~46 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~73 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[23]~46_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[23]~42_combout ),
	.cin(gnd),
	.combout(\pc_cntr~73_combout ),
	.cout());
defparam \pc_cntr~73 .lut_mask = 16'h5E0E;
defparam \pc_cntr~73 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~74 (
	.dataa(\mem_alu_out[23]~q ),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~73_combout ),
	.datad(\csr|mepc[23]~q ),
	.cin(gnd),
	.combout(\pc_cntr~74_combout ),
	.cout());
defparam \pc_cntr~74 .lut_mask = 16'hF838;
defparam \pc_cntr~74 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~75 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~74_combout ),
	.datac(\csr|mtvec[23]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~75_combout ),
	.cout());
defparam \pc_cntr~75 .lut_mask = 16'h88A0;
defparam \pc_cntr~75 .sum_lutc_input = "datac";

dffeas \pc_cntr[23] (
	.clk(clk_clk),
	.d(\pc_cntr~75_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[23]~q ),
	.prn(vcc));
defparam \pc_cntr[23] .is_wysiwyg = "true";
defparam \pc_cntr[23] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~22 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[23]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~22_combout ),
	.cout());
defparam \id_pc~22 .lut_mask = 16'h8080;
defparam \id_pc~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~22 (
	.dataa(id_pc_24),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~22_combout ),
	.cout());
defparam \ex_pc~22 .lut_mask = 16'h8080;
defparam \ex_pc~22 .sum_lutc_input = "datac";

dffeas \ex_pc[24] (
	.clk(clk_clk),
	.d(\ex_pc~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[24]~q ),
	.prn(vcc));
defparam \ex_pc[24] .is_wysiwyg = "true";
defparam \ex_pc[24] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~22 (
	.dataa(\ex_pc[24]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~22_combout ),
	.cout());
defparam \mem_pc~22 .lut_mask = 16'h8888;
defparam \mem_pc~22 .sum_lutc_input = "datac";

dffeas \mem_pc[24] (
	.clk(clk_clk),
	.d(\mem_pc~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[24]~q ),
	.prn(vcc));
defparam \mem_pc[24] .is_wysiwyg = "true";
defparam \mem_pc[24] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~13 (
	.dataa(\ex_csr_addr[4]~q ),
	.datab(\ex_ctrl_imm_type.011~q ),
	.datac(\ex_csr_addr[11]~q ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\mem_imm~13_combout ),
	.cout());
defparam \mem_imm~13 .lut_mask = 16'h88B8;
defparam \mem_imm~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~39 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\mem_imm~13_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_imm~39_combout ),
	.cout());
defparam \mem_imm~39 .lut_mask = 16'h8888;
defparam \mem_imm~39 .sum_lutc_input = "datac";

dffeas \mem_imm[24] (
	.clk(clk_clk),
	.d(\mem_imm~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[24]~q ),
	.prn(vcc));
defparam \mem_imm[24] .is_wysiwyg = "true";
defparam \mem_imm[24] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[24]~48 (
	.dataa(\mem_pc[24]~q ),
	.datab(\mem_imm[24]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[23]~47 ),
	.combout(\_T_3862[24]~48_combout ),
	.cout(\_T_3862[24]~49 ));
defparam \_T_3862[24]~48 .lut_mask = 16'h698E;
defparam \_T_3862[24]~48 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \mem_csr_data~34 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[24]~216_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~34_combout ),
	.cout());
defparam \mem_csr_data~34 .lut_mask = 16'h8888;
defparam \mem_csr_data~34 .sum_lutc_input = "datac";

dffeas \mem_csr_data[24] (
	.clk(clk_clk),
	.d(\mem_csr_data~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[24]~q ),
	.prn(vcc));
defparam \mem_csr_data[24] .is_wysiwyg = "true";
defparam \mem_csr_data[24] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~28 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[24]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~28_combout ),
	.cout());
defparam \wb_csr_data~28 .lut_mask = 16'h8888;
defparam \wb_csr_data~28 .sum_lutc_input = "datac";

dffeas \wb_csr_data[24] (
	.clk(clk_clk),
	.d(\wb_csr_data~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[24]~q ),
	.prn(vcc));
defparam \wb_csr_data[24] .is_wysiwyg = "true";
defparam \wb_csr_data[24] .power_up = "low";

cyclone10lp_lcell_comb \npc[24]~44 (
	.dataa(\pc_cntr[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[23]~43 ),
	.combout(\npc[24]~44_combout ),
	.cout(\npc[24]~45 ));
defparam \npc[24]~44 .lut_mask = 16'hA50A;
defparam \npc[24]~44 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~28 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[24]~44_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~28_combout ),
	.cout());
defparam \id_npc~28 .lut_mask = 16'h8080;
defparam \id_npc~28 .sum_lutc_input = "datac";

dffeas \id_npc[24] (
	.clk(clk_clk),
	.d(\id_npc~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[24]~q ),
	.prn(vcc));
defparam \id_npc[24] .is_wysiwyg = "true";
defparam \id_npc[24] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~28 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[24]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~28_combout ),
	.cout());
defparam \ex_npc~28 .lut_mask = 16'h8080;
defparam \ex_npc~28 .sum_lutc_input = "datac";

dffeas \ex_npc[24] (
	.clk(clk_clk),
	.d(\ex_npc~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[24]~q ),
	.prn(vcc));
defparam \ex_npc[24] .is_wysiwyg = "true";
defparam \ex_npc[24] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~26 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[24]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~26_combout ),
	.cout());
defparam \mem_npc~26 .lut_mask = 16'h8888;
defparam \mem_npc~26 .sum_lutc_input = "datac";

dffeas \mem_npc[24] (
	.clk(clk_clk),
	.d(\mem_npc~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[24]~q ),
	.prn(vcc));
defparam \mem_npc[24] .is_wysiwyg = "true";
defparam \mem_npc[24] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~26 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[24]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~26_combout ),
	.cout());
defparam \wb_npc~26 .lut_mask = 16'h8888;
defparam \wb_npc~26 .sum_lutc_input = "datac";

dffeas \wb_npc[24] (
	.clk(clk_clk),
	.d(\wb_npc~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[24]~q ),
	.prn(vcc));
defparam \wb_npc[24] .is_wysiwyg = "true";
defparam \wb_npc[24] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~28 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[24]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~28_combout ),
	.cout());
defparam \wb_alu_out~28 .lut_mask = 16'h8888;
defparam \wb_alu_out~28 .sum_lutc_input = "datac";

dffeas \wb_alu_out[24] (
	.clk(clk_clk),
	.d(\wb_alu_out~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[24]~q ),
	.prn(vcc));
defparam \wb_alu_out[24] .is_wysiwyg = "true";
defparam \wb_alu_out[24] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[24]~59 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[24]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[24]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[24]~59_combout ),
	.cout());
defparam \_T_3543__T_3854_data[24]~59 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[24]~59 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~85 (
	.dataa(\wb_dmem_read_data~30_combout ),
	.datab(av_readdata_pre_24),
	.datac(\wb_dmem_read_data~23_combout ),
	.datad(\wb_dmem_read_data[22]~32_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~85_combout ),
	.cout());
defparam \wb_dmem_read_data~85 .lut_mask = 16'h00AE;
defparam \wb_dmem_read_data~85 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[24] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~85_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[24]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[24] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[24] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[24]~60 (
	.dataa(\wb_csr_data[24]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[24]~59_combout ),
	.datad(\wb_dmem_read_data[24]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[24]~60_combout ),
	.cout());
defparam \_T_3543__T_3854_data[24]~60 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[24]~60 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a8 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[24]~60_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_a_first_bit_number = 8;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_b_first_bit_number = 8;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a8 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~31 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a8~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~31_combout ),
	.cout());
defparam \ex_rs_1~31 .lut_mask = 16'h8888;
defparam \ex_rs_1~31 .sum_lutc_input = "datac";

dffeas \ex_rs_1[24] (
	.clk(clk_clk),
	.d(\ex_rs_1~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[24]~q ),
	.prn(vcc));
defparam \ex_rs_1[24] .is_wysiwyg = "true";
defparam \ex_rs_1[24] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[24]~112 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_24),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[24]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[24]~112_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[24]~112 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[24]~112 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[24]~113 (
	.dataa(\ex_rs_1[24]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[24]~112_combout ),
	.datad(\wb_csr_data[24]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[24]~113_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[24]~113 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[24]~113 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[24]~114 (
	.dataa(\mem_alu_out[24]~q ),
	.datab(\ex_reg_rs2_bypass[24]~113_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[24]~114_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[24]~114 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[24]~114 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[24]~115 (
	.dataa(\ex_reg_rs2_bypass[24]~114_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[24]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[24]~115_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[24]~115 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[24]~115 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[24]~88 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_reg_rs2_bypass[24]~115_combout ),
	.datad(\mem_imm~13_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[24]~88_combout ),
	.cout());
defparam \alu_io_op2[24]~88 .lut_mask = 16'hB380;
defparam \alu_io_op2[24]~88 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a8 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[24]~60_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a8_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_a_first_bit_number = 8;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_b_first_bit_number = 8;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a8 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~30 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a8~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~30_combout ),
	.cout());
defparam \ex_rs_0~30 .lut_mask = 16'h0080;
defparam \ex_rs_0~30 .sum_lutc_input = "datac";

dffeas \ex_rs_0[24] (
	.clk(clk_clk),
	.d(\ex_rs_0~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[24]~q ),
	.prn(vcc));
defparam \ex_rs_0[24] .is_wysiwyg = "true";
defparam \ex_rs_0[24] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[24]~122 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(av_readdata_pre_24),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\wb_alu_out[24]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[24]~122_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[24]~122 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[24]~122 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[24]~123 (
	.dataa(\ex_rs_0[24]~q ),
	.datab(\ex_reg_rs1_bypass[2]~138_combout ),
	.datac(\ex_reg_rs1_bypass[24]~122_combout ),
	.datad(\wb_csr_data[24]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[24]~123_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[24]~123 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[24]~123 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[24]~124 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[24]~123_combout ),
	.datad(\mem_csr_data[24]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[24]~124_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[24]~124 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[24]~124 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[24]~125 (
	.dataa(\ex_reg_rs1_bypass[24]~124_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[24]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[24]~125_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[24]~125 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[24]~125 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[24]~115 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[24]~q ),
	.datad(\ex_reg_rs1_bypass[24]~125_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[24]~115_combout ),
	.cout());
defparam \alu_io_op1[24]~115 .lut_mask = 16'h6240;
defparam \alu_io_op1[24]~115 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~133 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\alu_io_op2[24]~88_combout ),
	.datad(\alu_io_op1[24]~115_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~133_combout ),
	.cout());
defparam \mem_alu_out~133 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~133 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~134 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~133_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~240_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~134_combout ),
	.cout());
defparam \mem_alu_out~134 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~134 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~115 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[24]~115_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~134_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~115_combout ),
	.cout());
defparam \mem_alu_out~115 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~115 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~116 (
	.dataa(\alu_io_op2[24]~88_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~115_combout ),
	.datad(\alu|ShiftRight0~256_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~116_combout ),
	.cout());
defparam \mem_alu_out~116 .lut_mask = 16'hF838;
defparam \mem_alu_out~116 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~117 (
	.dataa(\mem_alu_out~116_combout ),
	.datab(\alu|_T_3[24]~48_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~117_combout ),
	.cout());
defparam \mem_alu_out~117 .lut_mask = 16'h00AC;
defparam \mem_alu_out~117 .sum_lutc_input = "datac";

dffeas \mem_alu_out[24] (
	.clk(clk_clk),
	.d(\mem_alu_out~117_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[24]~q ),
	.prn(vcc));
defparam \mem_alu_out[24] .is_wysiwyg = "true";
defparam \mem_alu_out[24] .power_up = "low";

cyclone10lp_lcell_comb \pc_cntr~76 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(\mem_alu_out[24]~q ),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[24]~44_combout ),
	.cin(gnd),
	.combout(\pc_cntr~76_combout ),
	.cout());
defparam \pc_cntr~76 .lut_mask = 16'hDAD0;
defparam \pc_cntr~76 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~77 (
	.dataa(\_T_3862[24]~48_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~76_combout ),
	.datad(\csr|mepc[24]~q ),
	.cin(gnd),
	.combout(\pc_cntr~77_combout ),
	.cout());
defparam \pc_cntr~77 .lut_mask = 16'hF2C2;
defparam \pc_cntr~77 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~78 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~77_combout ),
	.datac(\csr|mtvec[24]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~78_combout ),
	.cout());
defparam \pc_cntr~78 .lut_mask = 16'h88A0;
defparam \pc_cntr~78 .sum_lutc_input = "datac";

dffeas \pc_cntr[24] (
	.clk(clk_clk),
	.d(\pc_cntr~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[24]~q ),
	.prn(vcc));
defparam \pc_cntr[24] .is_wysiwyg = "true";
defparam \pc_cntr[24] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~23 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[24]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~23_combout ),
	.cout());
defparam \id_pc~23 .lut_mask = 16'h8080;
defparam \id_pc~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~23 (
	.dataa(id_pc_25),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~23_combout ),
	.cout());
defparam \ex_pc~23 .lut_mask = 16'h8080;
defparam \ex_pc~23 .sum_lutc_input = "datac";

dffeas \ex_pc[25] (
	.clk(clk_clk),
	.d(\ex_pc~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[25]~q ),
	.prn(vcc));
defparam \ex_pc[25] .is_wysiwyg = "true";
defparam \ex_pc[25] .power_up = "low";

cyclone10lp_lcell_comb \npc[25]~46 (
	.dataa(\pc_cntr[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[24]~45 ),
	.combout(\npc[25]~46_combout ),
	.cout(\npc[25]~47 ));
defparam \npc[25]~46 .lut_mask = 16'h5A5F;
defparam \npc[25]~46 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~29 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[25]~46_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~29_combout ),
	.cout());
defparam \id_npc~29 .lut_mask = 16'h8080;
defparam \id_npc~29 .sum_lutc_input = "datac";

dffeas \id_npc[25] (
	.clk(clk_clk),
	.d(\id_npc~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[25]~q ),
	.prn(vcc));
defparam \id_npc[25] .is_wysiwyg = "true";
defparam \id_npc[25] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~29 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[25]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~29_combout ),
	.cout());
defparam \ex_npc~29 .lut_mask = 16'h8080;
defparam \ex_npc~29 .sum_lutc_input = "datac";

dffeas \ex_npc[25] (
	.clk(clk_clk),
	.d(\ex_npc~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[25]~q ),
	.prn(vcc));
defparam \ex_npc[25] .is_wysiwyg = "true";
defparam \ex_npc[25] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~27 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[25]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~27_combout ),
	.cout());
defparam \mem_npc~27 .lut_mask = 16'h8888;
defparam \mem_npc~27 .sum_lutc_input = "datac";

dffeas \mem_npc[25] (
	.clk(clk_clk),
	.d(\mem_npc~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[25]~q ),
	.prn(vcc));
defparam \mem_npc[25] .is_wysiwyg = "true";
defparam \mem_npc[25] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~27 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[25]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~27_combout ),
	.cout());
defparam \wb_npc~27 .lut_mask = 16'h8888;
defparam \wb_npc~27 .sum_lutc_input = "datac";

dffeas \wb_npc[25] (
	.clk(clk_clk),
	.d(\wb_npc~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[25]~q ),
	.prn(vcc));
defparam \wb_npc[25] .is_wysiwyg = "true";
defparam \wb_npc[25] .power_up = "low";

cyclone10lp_lcell_comb \mem_csr_data~38 (
	.dataa(\csr|io_out[25]~221_combout ),
	.datab(\csr|io_out[25]~222_combout ),
	.datac(\mem_ctrl_mem_wr~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~38_combout ),
	.cout());
defparam \mem_csr_data~38 .lut_mask = 16'hE0E0;
defparam \mem_csr_data~38 .sum_lutc_input = "datac";

dffeas \mem_csr_data[25] (
	.clk(clk_clk),
	.d(\mem_csr_data~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[25]~q ),
	.prn(vcc));
defparam \mem_csr_data[25] .is_wysiwyg = "true";
defparam \mem_csr_data[25] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~29 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[25]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~29_combout ),
	.cout());
defparam \wb_csr_data~29 .lut_mask = 16'h8888;
defparam \wb_csr_data~29 .sum_lutc_input = "datac";

dffeas \wb_csr_data[25] (
	.clk(clk_clk),
	.d(\wb_csr_data~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[25]~q ),
	.prn(vcc));
defparam \wb_csr_data[25] .is_wysiwyg = "true";
defparam \wb_csr_data[25] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~29 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[25]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~29_combout ),
	.cout());
defparam \wb_alu_out~29 .lut_mask = 16'h8888;
defparam \wb_alu_out~29 .sum_lutc_input = "datac";

dffeas \wb_alu_out[25] (
	.clk(clk_clk),
	.d(\wb_alu_out~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[25]~q ),
	.prn(vcc));
defparam \wb_alu_out[25] .is_wysiwyg = "true";
defparam \wb_alu_out[25] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[25]~61 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[25]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[25]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[25]~61_combout ),
	.cout());
defparam \_T_3543__T_3854_data[25]~61 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[25]~61 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~86 (
	.dataa(\wb_dmem_read_data~36_combout ),
	.datab(av_readdata_pre_25),
	.datac(\wb_dmem_read_data~23_combout ),
	.datad(\wb_dmem_read_data[22]~32_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~86_combout ),
	.cout());
defparam \wb_dmem_read_data~86 .lut_mask = 16'h00AE;
defparam \wb_dmem_read_data~86 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[25] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~86_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[25]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[25] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[25] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[25]~62 (
	.dataa(\wb_npc[25]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[25]~61_combout ),
	.datad(\wb_dmem_read_data[25]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[25]~62_combout ),
	.cout());
defparam \_T_3543__T_3854_data[25]~62 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[25]~62 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a7 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[25]~62_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a7_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_a_first_bit_number = 7;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_b_first_bit_number = 7;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a7 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~31 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a7~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~31_combout ),
	.cout());
defparam \ex_rs_0~31 .lut_mask = 16'h0080;
defparam \ex_rs_0~31 .sum_lutc_input = "datac";

dffeas \ex_rs_0[25] (
	.clk(clk_clk),
	.d(\ex_rs_0~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[25]~q ),
	.prn(vcc));
defparam \ex_rs_0[25] .is_wysiwyg = "true";
defparam \ex_rs_0[25] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[25]~126 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(\ex_rs_0[25]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\wb_alu_out[25]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[25]~126_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[25]~126 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[25]~126 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[25]~127 (
	.dataa(av_readdata_pre_25),
	.datab(\ex_reg_rs1_bypass[2]~7_combout ),
	.datac(\ex_reg_rs1_bypass[25]~126_combout ),
	.datad(\wb_csr_data[25]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[25]~127_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[25]~127 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[25]~127 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[25]~128 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[25]~127_combout ),
	.datad(\mem_csr_data[25]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[25]~128_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[25]~128 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[25]~128 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[25]~129 (
	.dataa(\ex_reg_rs1_bypass[25]~128_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[25]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[25]~129_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[25]~129 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[25]~129 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[25]~116 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[25]~q ),
	.datad(\ex_reg_rs1_bypass[25]~129_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[25]~116_combout ),
	.cout());
defparam \alu_io_op1[25]~116 .lut_mask = 16'h6240;
defparam \alu_io_op1[25]~116 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a7 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[25]~62_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_a_first_bit_number = 7;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_b_first_bit_number = 7;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a7 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~30 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a7~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~30_combout ),
	.cout());
defparam \ex_rs_1~30 .lut_mask = 16'h8888;
defparam \ex_rs_1~30 .sum_lutc_input = "datac";

dffeas \ex_rs_1[25] (
	.clk(clk_clk),
	.d(\ex_rs_1~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[25]~q ),
	.prn(vcc));
defparam \ex_rs_1[25] .is_wysiwyg = "true";
defparam \ex_rs_1[25] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[25]~108 (
	.dataa(\ex_reg_rs2_bypass[7]~5_combout ),
	.datab(\ex_rs_1[25]~q ),
	.datac(\ex_reg_rs2_bypass[7]~4_combout ),
	.datad(\wb_alu_out[25]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[25]~108_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[25]~108 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[25]~108 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[25]~109 (
	.dataa(av_readdata_pre_25),
	.datab(\ex_reg_rs2_bypass[7]~5_combout ),
	.datac(\ex_reg_rs2_bypass[25]~108_combout ),
	.datad(\wb_csr_data[25]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[25]~109_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[25]~109 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[25]~109 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[25]~110 (
	.dataa(\mem_alu_out[25]~q ),
	.datab(\ex_reg_rs2_bypass[25]~109_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[25]~110_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[25]~110 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[25]~110 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[25]~111 (
	.dataa(\ex_reg_rs2_bypass[25]~110_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[25]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[25]~111_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[25]~111 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[25]~111 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~12 (
	.dataa(\ex_csr_addr[5]~q ),
	.datab(\ex_ctrl_imm_type.011~q ),
	.datac(\ex_csr_addr[11]~q ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\mem_imm~12_combout ),
	.cout());
defparam \mem_imm~12 .lut_mask = 16'h88B8;
defparam \mem_imm~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[25]~87 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_reg_rs2_bypass[25]~111_combout ),
	.datad(\mem_imm~12_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[25]~87_combout ),
	.cout());
defparam \alu_io_op2[25]~87 .lut_mask = 16'hB380;
defparam \alu_io_op2[25]~87 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~118 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\alu|_T_123[25]~combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~236_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~118_combout ),
	.cout());
defparam \mem_alu_out~118 .lut_mask = 16'hDAD0;
defparam \mem_alu_out~118 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~119 (
	.dataa(\alu_io_op1[25]~116_combout ),
	.datab(\alu_io_op2[25]~87_combout ),
	.datac(\mem_alu_out~118_combout ),
	.datad(\alu|LessThan0~0_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~119_combout ),
	.cout());
defparam \mem_alu_out~119 .lut_mask = 16'hF08E;
defparam \mem_alu_out~119 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~120 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[25]~87_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~119_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~120_combout ),
	.cout());
defparam \mem_alu_out~120 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~120 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~121 (
	.dataa(\alu_io_op1[25]~116_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~120_combout ),
	.datad(\alu|ShiftRight0~254_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~121_combout ),
	.cout());
defparam \mem_alu_out~121 .lut_mask = 16'hF838;
defparam \mem_alu_out~121 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~122 (
	.dataa(\mem_alu_out~121_combout ),
	.datab(\alu|_T_3[25]~50_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~122_combout ),
	.cout());
defparam \mem_alu_out~122 .lut_mask = 16'h00AC;
defparam \mem_alu_out~122 .sum_lutc_input = "datac";

dffeas \mem_alu_out[25] (
	.clk(clk_clk),
	.d(\mem_alu_out~122_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[25]~q ),
	.prn(vcc));
defparam \mem_alu_out[25] .is_wysiwyg = "true";
defparam \mem_alu_out[25] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~23 (
	.dataa(\ex_pc[25]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~23_combout ),
	.cout());
defparam \mem_pc~23 .lut_mask = 16'h8888;
defparam \mem_pc~23 .sum_lutc_input = "datac";

dffeas \mem_pc[25] (
	.clk(clk_clk),
	.d(\mem_pc~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[25]~q ),
	.prn(vcc));
defparam \mem_pc[25] .is_wysiwyg = "true";
defparam \mem_pc[25] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~40 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\mem_imm~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_imm~40_combout ),
	.cout());
defparam \mem_imm~40 .lut_mask = 16'h8888;
defparam \mem_imm~40 .sum_lutc_input = "datac";

dffeas \mem_imm[25] (
	.clk(clk_clk),
	.d(\mem_imm~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[25]~q ),
	.prn(vcc));
defparam \mem_imm[25] .is_wysiwyg = "true";
defparam \mem_imm[25] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[25]~50 (
	.dataa(\mem_pc[25]~q ),
	.datab(\mem_imm[25]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[24]~49 ),
	.combout(\_T_3862[25]~50_combout ),
	.cout(\_T_3862[25]~51 ));
defparam \_T_3862[25]~50 .lut_mask = 16'h9617;
defparam \_T_3862[25]~50 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~79 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[25]~50_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[25]~46_combout ),
	.cin(gnd),
	.combout(\pc_cntr~79_combout ),
	.cout());
defparam \pc_cntr~79 .lut_mask = 16'h5E0E;
defparam \pc_cntr~79 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~80 (
	.dataa(\mem_alu_out[25]~q ),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~79_combout ),
	.datad(\csr|mepc[25]~q ),
	.cin(gnd),
	.combout(\pc_cntr~80_combout ),
	.cout());
defparam \pc_cntr~80 .lut_mask = 16'hF838;
defparam \pc_cntr~80 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~81 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~80_combout ),
	.datac(\csr|mtvec[25]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~81_combout ),
	.cout());
defparam \pc_cntr~81 .lut_mask = 16'h88A0;
defparam \pc_cntr~81 .sum_lutc_input = "datac";

dffeas \pc_cntr[25] (
	.clk(clk_clk),
	.d(\pc_cntr~81_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[25]~q ),
	.prn(vcc));
defparam \pc_cntr[25] .is_wysiwyg = "true";
defparam \pc_cntr[25] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~24 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[25]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~24_combout ),
	.cout());
defparam \id_pc~24 .lut_mask = 16'h8080;
defparam \id_pc~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~24 (
	.dataa(id_pc_26),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~24_combout ),
	.cout());
defparam \ex_pc~24 .lut_mask = 16'h8080;
defparam \ex_pc~24 .sum_lutc_input = "datac";

dffeas \ex_pc[26] (
	.clk(clk_clk),
	.d(\ex_pc~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[26]~q ),
	.prn(vcc));
defparam \ex_pc[26] .is_wysiwyg = "true";
defparam \ex_pc[26] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~24 (
	.dataa(\ex_pc[26]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~24_combout ),
	.cout());
defparam \mem_pc~24 .lut_mask = 16'h8888;
defparam \mem_pc~24 .sum_lutc_input = "datac";

dffeas \mem_pc[26] (
	.clk(clk_clk),
	.d(\mem_pc~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[26]~q ),
	.prn(vcc));
defparam \mem_pc[26] .is_wysiwyg = "true";
defparam \mem_pc[26] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~14 (
	.dataa(\ex_csr_addr[6]~q ),
	.datab(\ex_ctrl_imm_type.011~q ),
	.datac(\ex_csr_addr[11]~q ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\mem_imm~14_combout ),
	.cout());
defparam \mem_imm~14 .lut_mask = 16'h88B8;
defparam \mem_imm~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~41 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\mem_imm~14_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_imm~41_combout ),
	.cout());
defparam \mem_imm~41 .lut_mask = 16'h8888;
defparam \mem_imm~41 .sum_lutc_input = "datac";

dffeas \mem_imm[26] (
	.clk(clk_clk),
	.d(\mem_imm~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[26]~q ),
	.prn(vcc));
defparam \mem_imm[26] .is_wysiwyg = "true";
defparam \mem_imm[26] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[26]~52 (
	.dataa(\mem_pc[26]~q ),
	.datab(\mem_imm[26]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[25]~51 ),
	.combout(\_T_3862[26]~52_combout ),
	.cout(\_T_3862[26]~53 ));
defparam \_T_3862[26]~52 .lut_mask = 16'h698E;
defparam \_T_3862[26]~52 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \mem_csr_data~35 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[26]~230_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~35_combout ),
	.cout());
defparam \mem_csr_data~35 .lut_mask = 16'h8888;
defparam \mem_csr_data~35 .sum_lutc_input = "datac";

dffeas \mem_csr_data[26] (
	.clk(clk_clk),
	.d(\mem_csr_data~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[26]~q ),
	.prn(vcc));
defparam \mem_csr_data[26] .is_wysiwyg = "true";
defparam \mem_csr_data[26] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~30 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[26]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~30_combout ),
	.cout());
defparam \wb_csr_data~30 .lut_mask = 16'h8888;
defparam \wb_csr_data~30 .sum_lutc_input = "datac";

dffeas \wb_csr_data[26] (
	.clk(clk_clk),
	.d(\wb_csr_data~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[26]~q ),
	.prn(vcc));
defparam \wb_csr_data[26] .is_wysiwyg = "true";
defparam \wb_csr_data[26] .power_up = "low";

cyclone10lp_lcell_comb \npc[26]~48 (
	.dataa(\pc_cntr[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[25]~47 ),
	.combout(\npc[26]~48_combout ),
	.cout(\npc[26]~49 ));
defparam \npc[26]~48 .lut_mask = 16'hA50A;
defparam \npc[26]~48 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~30 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[26]~48_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~30_combout ),
	.cout());
defparam \id_npc~30 .lut_mask = 16'h8080;
defparam \id_npc~30 .sum_lutc_input = "datac";

dffeas \id_npc[26] (
	.clk(clk_clk),
	.d(\id_npc~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[26]~q ),
	.prn(vcc));
defparam \id_npc[26] .is_wysiwyg = "true";
defparam \id_npc[26] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~30 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[26]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~30_combout ),
	.cout());
defparam \ex_npc~30 .lut_mask = 16'h8080;
defparam \ex_npc~30 .sum_lutc_input = "datac";

dffeas \ex_npc[26] (
	.clk(clk_clk),
	.d(\ex_npc~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[26]~q ),
	.prn(vcc));
defparam \ex_npc[26] .is_wysiwyg = "true";
defparam \ex_npc[26] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~28 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[26]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~28_combout ),
	.cout());
defparam \mem_npc~28 .lut_mask = 16'h8888;
defparam \mem_npc~28 .sum_lutc_input = "datac";

dffeas \mem_npc[26] (
	.clk(clk_clk),
	.d(\mem_npc~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[26]~q ),
	.prn(vcc));
defparam \mem_npc[26] .is_wysiwyg = "true";
defparam \mem_npc[26] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~28 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[26]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~28_combout ),
	.cout());
defparam \wb_npc~28 .lut_mask = 16'h8888;
defparam \wb_npc~28 .sum_lutc_input = "datac";

dffeas \wb_npc[26] (
	.clk(clk_clk),
	.d(\wb_npc~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[26]~q ),
	.prn(vcc));
defparam \wb_npc[26] .is_wysiwyg = "true";
defparam \wb_npc[26] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~30 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[26]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~30_combout ),
	.cout());
defparam \wb_alu_out~30 .lut_mask = 16'h8888;
defparam \wb_alu_out~30 .sum_lutc_input = "datac";

dffeas \wb_alu_out[26] (
	.clk(clk_clk),
	.d(\wb_alu_out~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[26]~q ),
	.prn(vcc));
defparam \wb_alu_out[26] .is_wysiwyg = "true";
defparam \wb_alu_out[26] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[26]~63 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[26]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[26]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[26]~63_combout ),
	.cout());
defparam \_T_3543__T_3854_data[26]~63 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[26]~63 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~87 (
	.dataa(\wb_dmem_read_data~30_combout ),
	.datab(av_readdata_pre_26),
	.datac(\wb_dmem_read_data~23_combout ),
	.datad(\wb_dmem_read_data[22]~32_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~87_combout ),
	.cout());
defparam \wb_dmem_read_data~87 .lut_mask = 16'h00AE;
defparam \wb_dmem_read_data~87 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[26] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~87_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[26]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[26] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[26] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[26]~64 (
	.dataa(\wb_csr_data[26]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[26]~63_combout ),
	.datad(\wb_dmem_read_data[26]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[26]~64_combout ),
	.cout());
defparam \_T_3543__T_3854_data[26]~64 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[26]~64 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a6 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[26]~64_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_a_first_bit_number = 6;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_b_first_bit_number = 6;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a6 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~32 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a6~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~32_combout ),
	.cout());
defparam \ex_rs_1~32 .lut_mask = 16'h8888;
defparam \ex_rs_1~32 .sum_lutc_input = "datac";

dffeas \ex_rs_1[26] (
	.clk(clk_clk),
	.d(\ex_rs_1~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[26]~q ),
	.prn(vcc));
defparam \ex_rs_1[26] .is_wysiwyg = "true";
defparam \ex_rs_1[26] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[26]~116 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_26),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[26]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[26]~116_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[26]~116 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[26]~116 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[26]~117 (
	.dataa(\ex_rs_1[26]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[26]~116_combout ),
	.datad(\wb_csr_data[26]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[26]~117_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[26]~117 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[26]~117 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[26]~118 (
	.dataa(\mem_alu_out[26]~q ),
	.datab(\ex_reg_rs2_bypass[26]~117_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[26]~118_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[26]~118 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[26]~118 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[26]~119 (
	.dataa(\ex_reg_rs2_bypass[26]~118_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[26]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[26]~119_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[26]~119 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[26]~119 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[26]~89 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_reg_rs2_bypass[26]~119_combout ),
	.datad(\mem_imm~14_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[26]~89_combout ),
	.cout());
defparam \alu_io_op2[26]~89 .lut_mask = 16'hB380;
defparam \alu_io_op2[26]~89 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a6 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[26]~64_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a6_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_a_first_bit_number = 6;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_b_first_bit_number = 6;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a6 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~32 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a6~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~32_combout ),
	.cout());
defparam \ex_rs_0~32 .lut_mask = 16'h0080;
defparam \ex_rs_0~32 .sum_lutc_input = "datac";

dffeas \ex_rs_0[26] (
	.clk(clk_clk),
	.d(\ex_rs_0~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[26]~q ),
	.prn(vcc));
defparam \ex_rs_0[26] .is_wysiwyg = "true";
defparam \ex_rs_0[26] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[26]~130 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(av_readdata_pre_26),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\wb_alu_out[26]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[26]~130_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[26]~130 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[26]~130 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[26]~131 (
	.dataa(\ex_rs_0[26]~q ),
	.datab(\ex_reg_rs1_bypass[2]~138_combout ),
	.datac(\ex_reg_rs1_bypass[26]~130_combout ),
	.datad(\wb_csr_data[26]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[26]~131_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[26]~131 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[26]~131 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[26]~132 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[26]~131_combout ),
	.datad(\mem_csr_data[26]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[26]~132_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[26]~132 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[26]~132 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[26]~133 (
	.dataa(\ex_reg_rs1_bypass[26]~132_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[26]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[26]~133_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[26]~133 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[26]~133 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[26]~117 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[26]~q ),
	.datad(\ex_reg_rs1_bypass[26]~133_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[26]~117_combout ),
	.cout());
defparam \alu_io_op1[26]~117 .lut_mask = 16'h6240;
defparam \alu_io_op1[26]~117 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~131 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\alu_io_op2[26]~89_combout ),
	.datad(\alu_io_op1[26]~117_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~131_combout ),
	.cout());
defparam \mem_alu_out~131 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~131 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~132 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~131_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~233_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~132_combout ),
	.cout());
defparam \mem_alu_out~132 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~132 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~123 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[26]~117_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~132_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~123_combout ),
	.cout());
defparam \mem_alu_out~123 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~123 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~124 (
	.dataa(\alu_io_op2[26]~89_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~123_combout ),
	.datad(\alu|ShiftRight0~253_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~124_combout ),
	.cout());
defparam \mem_alu_out~124 .lut_mask = 16'hF838;
defparam \mem_alu_out~124 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~125 (
	.dataa(\mem_alu_out~124_combout ),
	.datab(\alu|_T_3[26]~52_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~125_combout ),
	.cout());
defparam \mem_alu_out~125 .lut_mask = 16'h00AC;
defparam \mem_alu_out~125 .sum_lutc_input = "datac";

dffeas \mem_alu_out[26] (
	.clk(clk_clk),
	.d(\mem_alu_out~125_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[26]~q ),
	.prn(vcc));
defparam \mem_alu_out[26] .is_wysiwyg = "true";
defparam \mem_alu_out[26] .power_up = "low";

cyclone10lp_lcell_comb \pc_cntr~82 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(\mem_alu_out[26]~q ),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[26]~48_combout ),
	.cin(gnd),
	.combout(\pc_cntr~82_combout ),
	.cout());
defparam \pc_cntr~82 .lut_mask = 16'hDAD0;
defparam \pc_cntr~82 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~83 (
	.dataa(\_T_3862[26]~52_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~82_combout ),
	.datad(\csr|mepc[26]~q ),
	.cin(gnd),
	.combout(\pc_cntr~83_combout ),
	.cout());
defparam \pc_cntr~83 .lut_mask = 16'hF2C2;
defparam \pc_cntr~83 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~84 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~83_combout ),
	.datac(\csr|mtvec[26]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~84_combout ),
	.cout());
defparam \pc_cntr~84 .lut_mask = 16'h88A0;
defparam \pc_cntr~84 .sum_lutc_input = "datac";

dffeas \pc_cntr[26] (
	.clk(clk_clk),
	.d(\pc_cntr~84_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[26]~q ),
	.prn(vcc));
defparam \pc_cntr[26] .is_wysiwyg = "true";
defparam \pc_cntr[26] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~25 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[26]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~25_combout ),
	.cout());
defparam \id_pc~25 .lut_mask = 16'h8080;
defparam \id_pc~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~25 (
	.dataa(id_pc_27),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~25_combout ),
	.cout());
defparam \ex_pc~25 .lut_mask = 16'h8080;
defparam \ex_pc~25 .sum_lutc_input = "datac";

dffeas \ex_pc[27] (
	.clk(clk_clk),
	.d(\ex_pc~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[27]~q ),
	.prn(vcc));
defparam \ex_pc[27] .is_wysiwyg = "true";
defparam \ex_pc[27] .power_up = "low";

cyclone10lp_lcell_comb \npc[27]~50 (
	.dataa(\pc_cntr[27]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[26]~49 ),
	.combout(\npc[27]~50_combout ),
	.cout(\npc[27]~51 ));
defparam \npc[27]~50 .lut_mask = 16'h5A5F;
defparam \npc[27]~50 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~31 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[27]~50_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~31_combout ),
	.cout());
defparam \id_npc~31 .lut_mask = 16'h8080;
defparam \id_npc~31 .sum_lutc_input = "datac";

dffeas \id_npc[27] (
	.clk(clk_clk),
	.d(\id_npc~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[27]~q ),
	.prn(vcc));
defparam \id_npc[27] .is_wysiwyg = "true";
defparam \id_npc[27] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~31 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[27]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~31_combout ),
	.cout());
defparam \ex_npc~31 .lut_mask = 16'h8080;
defparam \ex_npc~31 .sum_lutc_input = "datac";

dffeas \ex_npc[27] (
	.clk(clk_clk),
	.d(\ex_npc~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[27]~q ),
	.prn(vcc));
defparam \ex_npc[27] .is_wysiwyg = "true";
defparam \ex_npc[27] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~29 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[27]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~29_combout ),
	.cout());
defparam \mem_npc~29 .lut_mask = 16'h8888;
defparam \mem_npc~29 .sum_lutc_input = "datac";

dffeas \mem_npc[27] (
	.clk(clk_clk),
	.d(\mem_npc~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[27]~q ),
	.prn(vcc));
defparam \mem_npc[27] .is_wysiwyg = "true";
defparam \mem_npc[27] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~29 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[27]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~29_combout ),
	.cout());
defparam \wb_npc~29 .lut_mask = 16'h8888;
defparam \wb_npc~29 .sum_lutc_input = "datac";

dffeas \wb_npc[27] (
	.clk(clk_clk),
	.d(\wb_npc~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[27]~q ),
	.prn(vcc));
defparam \wb_npc[27] .is_wysiwyg = "true";
defparam \wb_npc[27] .power_up = "low";

cyclone10lp_lcell_comb \mem_csr_data~39 (
	.dataa(\csr|io_out[27]~235_combout ),
	.datab(\csr|io_out[27]~236_combout ),
	.datac(\mem_ctrl_mem_wr~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~39_combout ),
	.cout());
defparam \mem_csr_data~39 .lut_mask = 16'hE0E0;
defparam \mem_csr_data~39 .sum_lutc_input = "datac";

dffeas \mem_csr_data[27] (
	.clk(clk_clk),
	.d(\mem_csr_data~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[27]~q ),
	.prn(vcc));
defparam \mem_csr_data[27] .is_wysiwyg = "true";
defparam \mem_csr_data[27] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~31 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[27]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~31_combout ),
	.cout());
defparam \wb_csr_data~31 .lut_mask = 16'h8888;
defparam \wb_csr_data~31 .sum_lutc_input = "datac";

dffeas \wb_csr_data[27] (
	.clk(clk_clk),
	.d(\wb_csr_data~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[27]~q ),
	.prn(vcc));
defparam \wb_csr_data[27] .is_wysiwyg = "true";
defparam \wb_csr_data[27] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~31 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[27]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~31_combout ),
	.cout());
defparam \wb_alu_out~31 .lut_mask = 16'h8888;
defparam \wb_alu_out~31 .sum_lutc_input = "datac";

dffeas \wb_alu_out[27] (
	.clk(clk_clk),
	.d(\wb_alu_out~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[27]~q ),
	.prn(vcc));
defparam \wb_alu_out[27] .is_wysiwyg = "true";
defparam \wb_alu_out[27] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[27]~65 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[27]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[27]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[27]~65_combout ),
	.cout());
defparam \_T_3543__T_3854_data[27]~65 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[27]~65 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~88 (
	.dataa(\wb_dmem_read_data~36_combout ),
	.datab(av_readdata_pre_27),
	.datac(\wb_dmem_read_data~23_combout ),
	.datad(\wb_dmem_read_data[22]~32_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~88_combout ),
	.cout());
defparam \wb_dmem_read_data~88 .lut_mask = 16'h00AE;
defparam \wb_dmem_read_data~88 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[27] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~88_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[27]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[27] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[27] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[27]~66 (
	.dataa(\wb_npc[27]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[27]~65_combout ),
	.datad(\wb_dmem_read_data[27]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[27]~66_combout ),
	.cout());
defparam \_T_3543__T_3854_data[27]~66 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[27]~66 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a5 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[27]~66_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a5_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_a_first_bit_number = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_b_first_bit_number = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a5 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~33 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a5~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~33_combout ),
	.cout());
defparam \ex_rs_0~33 .lut_mask = 16'h0080;
defparam \ex_rs_0~33 .sum_lutc_input = "datac";

dffeas \ex_rs_0[27] (
	.clk(clk_clk),
	.d(\ex_rs_0~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[27]~q ),
	.prn(vcc));
defparam \ex_rs_0[27] .is_wysiwyg = "true";
defparam \ex_rs_0[27] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[27]~134 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(\ex_rs_0[27]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\wb_alu_out[27]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[27]~134_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[27]~134 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[27]~134 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[27]~135 (
	.dataa(av_readdata_pre_27),
	.datab(\ex_reg_rs1_bypass[2]~7_combout ),
	.datac(\ex_reg_rs1_bypass[27]~134_combout ),
	.datad(\wb_csr_data[27]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[27]~135_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[27]~135 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[27]~135 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[27]~136 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[27]~135_combout ),
	.datad(\mem_csr_data[27]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[27]~136_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[27]~136 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[27]~136 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[27]~137 (
	.dataa(\ex_reg_rs1_bypass[27]~136_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[27]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[27]~137_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[27]~137 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[27]~137 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[27]~118 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[27]~q ),
	.datad(\ex_reg_rs1_bypass[27]~137_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[27]~118_combout ),
	.cout());
defparam \alu_io_op1[27]~118 .lut_mask = 16'h6240;
defparam \alu_io_op1[27]~118 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a5 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[27]~66_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_a_first_bit_number = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_b_first_bit_number = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a5 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~33 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a5~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~33_combout ),
	.cout());
defparam \ex_rs_1~33 .lut_mask = 16'h8888;
defparam \ex_rs_1~33 .sum_lutc_input = "datac";

dffeas \ex_rs_1[27] (
	.clk(clk_clk),
	.d(\ex_rs_1~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[27]~q ),
	.prn(vcc));
defparam \ex_rs_1[27] .is_wysiwyg = "true";
defparam \ex_rs_1[27] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[27]~120 (
	.dataa(\ex_reg_rs2_bypass[7]~5_combout ),
	.datab(\ex_rs_1[27]~q ),
	.datac(\ex_reg_rs2_bypass[7]~4_combout ),
	.datad(\wb_alu_out[27]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[27]~120_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[27]~120 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[27]~120 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[27]~121 (
	.dataa(av_readdata_pre_27),
	.datab(\ex_reg_rs2_bypass[7]~5_combout ),
	.datac(\ex_reg_rs2_bypass[27]~120_combout ),
	.datad(\wb_csr_data[27]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[27]~121_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[27]~121 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[27]~121 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[27]~122 (
	.dataa(\mem_alu_out[27]~q ),
	.datab(\ex_reg_rs2_bypass[27]~121_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[27]~122_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[27]~122 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[27]~122 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[27]~123 (
	.dataa(\ex_reg_rs2_bypass[27]~122_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[27]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[27]~123_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[27]~123 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[27]~123 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~15 (
	.dataa(\ex_csr_addr[7]~q ),
	.datab(\ex_ctrl_imm_type.011~q ),
	.datac(\ex_csr_addr[11]~q ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\mem_imm~15_combout ),
	.cout());
defparam \mem_imm~15 .lut_mask = 16'h88B8;
defparam \mem_imm~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[27]~90 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_reg_rs2_bypass[27]~123_combout ),
	.datad(\mem_imm~15_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[27]~90_combout ),
	.cout());
defparam \alu_io_op2[27]~90 .lut_mask = 16'hB380;
defparam \alu_io_op2[27]~90 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~126 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\alu|_T_123[27]~combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~228_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~126_combout ),
	.cout());
defparam \mem_alu_out~126 .lut_mask = 16'hDAD0;
defparam \mem_alu_out~126 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~127 (
	.dataa(\alu_io_op1[27]~118_combout ),
	.datab(\alu_io_op2[27]~90_combout ),
	.datac(\mem_alu_out~126_combout ),
	.datad(\alu|LessThan0~0_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~127_combout ),
	.cout());
defparam \mem_alu_out~127 .lut_mask = 16'hF08E;
defparam \mem_alu_out~127 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~128 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[27]~90_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~127_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~128_combout ),
	.cout());
defparam \mem_alu_out~128 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~128 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~129 (
	.dataa(\alu_io_op1[27]~118_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~128_combout ),
	.datad(\alu|ShiftRight0~251_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~129_combout ),
	.cout());
defparam \mem_alu_out~129 .lut_mask = 16'hF838;
defparam \mem_alu_out~129 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~130 (
	.dataa(\mem_alu_out~129_combout ),
	.datab(\alu|_T_3[27]~54_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~130_combout ),
	.cout());
defparam \mem_alu_out~130 .lut_mask = 16'h00AC;
defparam \mem_alu_out~130 .sum_lutc_input = "datac";

dffeas \mem_alu_out[27] (
	.clk(clk_clk),
	.d(\mem_alu_out~130_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[27]~q ),
	.prn(vcc));
defparam \mem_alu_out[27] .is_wysiwyg = "true";
defparam \mem_alu_out[27] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~25 (
	.dataa(\ex_pc[27]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~25_combout ),
	.cout());
defparam \mem_pc~25 .lut_mask = 16'h8888;
defparam \mem_pc~25 .sum_lutc_input = "datac";

dffeas \mem_pc[27] (
	.clk(clk_clk),
	.d(\mem_pc~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[27]~q ),
	.prn(vcc));
defparam \mem_pc[27] .is_wysiwyg = "true";
defparam \mem_pc[27] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~42 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\mem_imm~15_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_imm~42_combout ),
	.cout());
defparam \mem_imm~42 .lut_mask = 16'h8888;
defparam \mem_imm~42 .sum_lutc_input = "datac";

dffeas \mem_imm[27] (
	.clk(clk_clk),
	.d(\mem_imm~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[27]~q ),
	.prn(vcc));
defparam \mem_imm[27] .is_wysiwyg = "true";
defparam \mem_imm[27] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[27]~54 (
	.dataa(\mem_pc[27]~q ),
	.datab(\mem_imm[27]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[26]~53 ),
	.combout(\_T_3862[27]~54_combout ),
	.cout(\_T_3862[27]~55 ));
defparam \_T_3862[27]~54 .lut_mask = 16'h9617;
defparam \_T_3862[27]~54 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~85 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[27]~54_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[27]~50_combout ),
	.cin(gnd),
	.combout(\pc_cntr~85_combout ),
	.cout());
defparam \pc_cntr~85 .lut_mask = 16'h5E0E;
defparam \pc_cntr~85 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~86 (
	.dataa(\mem_alu_out[27]~q ),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~85_combout ),
	.datad(\csr|mepc[27]~q ),
	.cin(gnd),
	.combout(\pc_cntr~86_combout ),
	.cout());
defparam \pc_cntr~86 .lut_mask = 16'hF838;
defparam \pc_cntr~86 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~87 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~86_combout ),
	.datac(\csr|mtvec[27]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~87_combout ),
	.cout());
defparam \pc_cntr~87 .lut_mask = 16'h88A0;
defparam \pc_cntr~87 .sum_lutc_input = "datac";

dffeas \pc_cntr[27] (
	.clk(clk_clk),
	.d(\pc_cntr~87_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[27]~q ),
	.prn(vcc));
defparam \pc_cntr[27] .is_wysiwyg = "true";
defparam \pc_cntr[27] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~26 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[27]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~26_combout ),
	.cout());
defparam \id_pc~26 .lut_mask = 16'h8080;
defparam \id_pc~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~26 (
	.dataa(id_pc_28),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~26_combout ),
	.cout());
defparam \ex_pc~26 .lut_mask = 16'h8080;
defparam \ex_pc~26 .sum_lutc_input = "datac";

dffeas \ex_pc[28] (
	.clk(clk_clk),
	.d(\ex_pc~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[28]~q ),
	.prn(vcc));
defparam \ex_pc[28] .is_wysiwyg = "true";
defparam \ex_pc[28] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~26 (
	.dataa(\ex_pc[28]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~26_combout ),
	.cout());
defparam \mem_pc~26 .lut_mask = 16'h8888;
defparam \mem_pc~26 .sum_lutc_input = "datac";

dffeas \mem_pc[28] (
	.clk(clk_clk),
	.d(\mem_pc~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[28]~q ),
	.prn(vcc));
defparam \mem_pc[28] .is_wysiwyg = "true";
defparam \mem_pc[28] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~5 (
	.dataa(\ex_csr_addr[8]~q ),
	.datab(\ex_ctrl_imm_type.011~q ),
	.datac(\ex_csr_addr[11]~q ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\mem_imm~5_combout ),
	.cout());
defparam \mem_imm~5 .lut_mask = 16'h88B8;
defparam \mem_imm~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~43 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\mem_imm~5_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_imm~43_combout ),
	.cout());
defparam \mem_imm~43 .lut_mask = 16'h8888;
defparam \mem_imm~43 .sum_lutc_input = "datac";

dffeas \mem_imm[28] (
	.clk(clk_clk),
	.d(\mem_imm~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[28]~q ),
	.prn(vcc));
defparam \mem_imm[28] .is_wysiwyg = "true";
defparam \mem_imm[28] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[28]~56 (
	.dataa(\mem_pc[28]~q ),
	.datab(\mem_imm[28]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[27]~55 ),
	.combout(\_T_3862[28]~56_combout ),
	.cout(\_T_3862[28]~57 ));
defparam \_T_3862[28]~56 .lut_mask = 16'h698E;
defparam \_T_3862[28]~56 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \mem_csr_data~10 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[28]~31_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~10_combout ),
	.cout());
defparam \mem_csr_data~10 .lut_mask = 16'h8888;
defparam \mem_csr_data~10 .sum_lutc_input = "datac";

dffeas \mem_csr_data[28] (
	.clk(clk_clk),
	.d(\mem_csr_data~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[28]~q ),
	.prn(vcc));
defparam \mem_csr_data[28] .is_wysiwyg = "true";
defparam \mem_csr_data[28] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[28]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~2_combout ),
	.cout());
defparam \wb_csr_data~2 .lut_mask = 16'h8888;
defparam \wb_csr_data~2 .sum_lutc_input = "datac";

dffeas \wb_csr_data[28] (
	.clk(clk_clk),
	.d(\wb_csr_data~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[28]~q ),
	.prn(vcc));
defparam \wb_csr_data[28] .is_wysiwyg = "true";
defparam \wb_csr_data[28] .power_up = "low";

cyclone10lp_lcell_comb \npc[28]~52 (
	.dataa(\pc_cntr[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[27]~51 ),
	.combout(\npc[28]~52_combout ),
	.cout(\npc[28]~53 ));
defparam \npc[28]~52 .lut_mask = 16'hA50A;
defparam \npc[28]~52 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~2 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[28]~52_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~2_combout ),
	.cout());
defparam \id_npc~2 .lut_mask = 16'h8080;
defparam \id_npc~2 .sum_lutc_input = "datac";

dffeas \id_npc[28] (
	.clk(clk_clk),
	.d(\id_npc~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[28]~q ),
	.prn(vcc));
defparam \id_npc[28] .is_wysiwyg = "true";
defparam \id_npc[28] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~2 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[28]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~2_combout ),
	.cout());
defparam \ex_npc~2 .lut_mask = 16'h8080;
defparam \ex_npc~2 .sum_lutc_input = "datac";

dffeas \ex_npc[28] (
	.clk(clk_clk),
	.d(\ex_npc~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[28]~q ),
	.prn(vcc));
defparam \ex_npc[28] .is_wysiwyg = "true";
defparam \ex_npc[28] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~0 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[28]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~0_combout ),
	.cout());
defparam \mem_npc~0 .lut_mask = 16'h8888;
defparam \mem_npc~0 .sum_lutc_input = "datac";

dffeas \mem_npc[28] (
	.clk(clk_clk),
	.d(\mem_npc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[28]~q ),
	.prn(vcc));
defparam \mem_npc[28] .is_wysiwyg = "true";
defparam \mem_npc[28] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[28]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~0_combout ),
	.cout());
defparam \wb_npc~0 .lut_mask = 16'h8888;
defparam \wb_npc~0 .sum_lutc_input = "datac";

dffeas \wb_npc[28] (
	.clk(clk_clk),
	.d(\wb_npc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[28]~q ),
	.prn(vcc));
defparam \wb_npc[28] .is_wysiwyg = "true";
defparam \wb_npc[28] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[28]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~2_combout ),
	.cout());
defparam \wb_alu_out~2 .lut_mask = 16'h8888;
defparam \wb_alu_out~2 .sum_lutc_input = "datac";

dffeas \wb_alu_out[28] (
	.clk(clk_clk),
	.d(\wb_alu_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[28]~q ),
	.prn(vcc));
defparam \wb_alu_out[28] .is_wysiwyg = "true";
defparam \wb_alu_out[28] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[28]~7 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[28]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[28]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[28]~7_combout ),
	.cout());
defparam \_T_3543__T_3854_data[28]~7 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[28]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~33 (
	.dataa(\wb_dmem_read_data~30_combout ),
	.datab(av_readdata_pre_28),
	.datac(\wb_dmem_read_data~23_combout ),
	.datad(\wb_dmem_read_data[22]~32_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~33_combout ),
	.cout());
defparam \wb_dmem_read_data~33 .lut_mask = 16'h00AE;
defparam \wb_dmem_read_data~33 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[28] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[28]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[28] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[28] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[28]~8 (
	.dataa(\wb_csr_data[28]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[28]~7_combout ),
	.datad(\wb_dmem_read_data[28]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[28]~8_combout ),
	.cout());
defparam \_T_3543__T_3854_data[28]~8 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[28]~8 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a4 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[28]~8_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_a_first_bit_number = 4;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_b_first_bit_number = 4;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a4 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~5 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a4~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~5_combout ),
	.cout());
defparam \ex_rs_1~5 .lut_mask = 16'h8888;
defparam \ex_rs_1~5 .sum_lutc_input = "datac";

dffeas \ex_rs_1[28] (
	.clk(clk_clk),
	.d(\ex_rs_1~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[28]~q ),
	.prn(vcc));
defparam \ex_rs_1[28] .is_wysiwyg = "true";
defparam \ex_rs_1[28] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[28]~19 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_28),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[28]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[28]~19_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[28]~19 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[28]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[28]~20 (
	.dataa(\ex_rs_1[28]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[28]~19_combout ),
	.datad(\wb_csr_data[28]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[28]~20_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[28]~20 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[28]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[28]~21 (
	.dataa(\mem_alu_out[28]~q ),
	.datab(\ex_reg_rs2_bypass[28]~20_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[28]~21_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[28]~21 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[28]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[28]~22 (
	.dataa(\ex_reg_rs2_bypass[28]~21_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[28]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[28]~22_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[28]~22 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[28]~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[28]~74 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_reg_rs2_bypass[28]~22_combout ),
	.datad(\mem_imm~5_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[28]~74_combout ),
	.cout());
defparam \alu_io_op2[28]~74 .lut_mask = 16'hB380;
defparam \alu_io_op2[28]~74 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a4 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[28]~8_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a4_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_a_first_bit_number = 4;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_b_first_bit_number = 4;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a4 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~4 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a4~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~4_combout ),
	.cout());
defparam \ex_rs_0~4 .lut_mask = 16'h0080;
defparam \ex_rs_0~4 .sum_lutc_input = "datac";

dffeas \ex_rs_0[28] (
	.clk(clk_clk),
	.d(\ex_rs_0~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[28]~q ),
	.prn(vcc));
defparam \ex_rs_0[28] .is_wysiwyg = "true";
defparam \ex_rs_0[28] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[28]~17 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(av_readdata_pre_28),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\wb_alu_out[28]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[28]~17_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[28]~17 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[28]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[28]~18 (
	.dataa(\ex_rs_0[28]~q ),
	.datab(\ex_reg_rs1_bypass[2]~138_combout ),
	.datac(\ex_reg_rs1_bypass[28]~17_combout ),
	.datad(\wb_csr_data[28]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[28]~18_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[28]~18 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[28]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[28]~19 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[28]~18_combout ),
	.datad(\mem_csr_data[28]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[28]~19_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[28]~19 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[28]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[28]~21 (
	.dataa(\ex_reg_rs1_bypass[28]~19_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[28]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[28]~21_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[28]~21 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[28]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[28]~90 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[28]~q ),
	.datad(\ex_reg_rs1_bypass[28]~21_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[28]~90_combout ),
	.cout());
defparam \alu_io_op1[28]~90 .lut_mask = 16'h6240;
defparam \alu_io_op1[28]~90 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~159 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\alu_io_op2[28]~74_combout ),
	.datad(\alu_io_op1[28]~90_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~159_combout ),
	.cout());
defparam \mem_alu_out~159 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~159 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~160 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~159_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~167_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~160_combout ),
	.cout());
defparam \mem_alu_out~160 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~160 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~21 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[28]~90_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~160_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~21_combout ),
	.cout());
defparam \mem_alu_out~21 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~22 (
	.dataa(\alu_io_op2[28]~74_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~21_combout ),
	.datad(\alu|ShiftRight0~152_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~22_combout ),
	.cout());
defparam \mem_alu_out~22 .lut_mask = 16'hF838;
defparam \mem_alu_out~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~23 (
	.dataa(\mem_alu_out~22_combout ),
	.datab(\alu|_T_3[28]~56_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~23_combout ),
	.cout());
defparam \mem_alu_out~23 .lut_mask = 16'h00AC;
defparam \mem_alu_out~23 .sum_lutc_input = "datac";

dffeas \mem_alu_out[28] (
	.clk(clk_clk),
	.d(\mem_alu_out~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[28]~q ),
	.prn(vcc));
defparam \mem_alu_out[28] .is_wysiwyg = "true";
defparam \mem_alu_out[28] .power_up = "low";

cyclone10lp_lcell_comb \pc_cntr~88 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(\mem_alu_out[28]~q ),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[28]~52_combout ),
	.cin(gnd),
	.combout(\pc_cntr~88_combout ),
	.cout());
defparam \pc_cntr~88 .lut_mask = 16'hDAD0;
defparam \pc_cntr~88 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~89 (
	.dataa(\_T_3862[28]~56_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~88_combout ),
	.datad(\csr|mepc[28]~q ),
	.cin(gnd),
	.combout(\pc_cntr~89_combout ),
	.cout());
defparam \pc_cntr~89 .lut_mask = 16'hF2C2;
defparam \pc_cntr~89 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~90 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~89_combout ),
	.datac(\csr|mtvec[28]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~90_combout ),
	.cout());
defparam \pc_cntr~90 .lut_mask = 16'h88A0;
defparam \pc_cntr~90 .sum_lutc_input = "datac";

dffeas \pc_cntr[28] (
	.clk(clk_clk),
	.d(\pc_cntr~90_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[28]~q ),
	.prn(vcc));
defparam \pc_cntr[28] .is_wysiwyg = "true";
defparam \pc_cntr[28] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~27 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[28]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~27_combout ),
	.cout());
defparam \id_pc~27 .lut_mask = 16'h8080;
defparam \id_pc~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~27 (
	.dataa(id_pc_29),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~27_combout ),
	.cout());
defparam \ex_pc~27 .lut_mask = 16'h8080;
defparam \ex_pc~27 .sum_lutc_input = "datac";

dffeas \ex_pc[29] (
	.clk(clk_clk),
	.d(\ex_pc~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[29]~q ),
	.prn(vcc));
defparam \ex_pc[29] .is_wysiwyg = "true";
defparam \ex_pc[29] .power_up = "low";

cyclone10lp_lcell_comb \npc[29]~54 (
	.dataa(\pc_cntr[29]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[28]~53 ),
	.combout(\npc[29]~54_combout ),
	.cout(\npc[29]~55 ));
defparam \npc[29]~54 .lut_mask = 16'h5A5F;
defparam \npc[29]~54 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~3 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[29]~54_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~3_combout ),
	.cout());
defparam \id_npc~3 .lut_mask = 16'h8080;
defparam \id_npc~3 .sum_lutc_input = "datac";

dffeas \id_npc[29] (
	.clk(clk_clk),
	.d(\id_npc~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[29]~q ),
	.prn(vcc));
defparam \id_npc[29] .is_wysiwyg = "true";
defparam \id_npc[29] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~3 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[29]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~3_combout ),
	.cout());
defparam \ex_npc~3 .lut_mask = 16'h8080;
defparam \ex_npc~3 .sum_lutc_input = "datac";

dffeas \ex_npc[29] (
	.clk(clk_clk),
	.d(\ex_npc~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[29]~q ),
	.prn(vcc));
defparam \ex_npc[29] .is_wysiwyg = "true";
defparam \ex_npc[29] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~1 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[29]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~1_combout ),
	.cout());
defparam \mem_npc~1 .lut_mask = 16'h8888;
defparam \mem_npc~1 .sum_lutc_input = "datac";

dffeas \mem_npc[29] (
	.clk(clk_clk),
	.d(\mem_npc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[29]~q ),
	.prn(vcc));
defparam \mem_npc[29] .is_wysiwyg = "true";
defparam \mem_npc[29] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~1 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[29]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~1_combout ),
	.cout());
defparam \wb_npc~1 .lut_mask = 16'h8888;
defparam \wb_npc~1 .sum_lutc_input = "datac";

dffeas \wb_npc[29] (
	.clk(clk_clk),
	.d(\wb_npc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[29]~q ),
	.prn(vcc));
defparam \wb_npc[29] .is_wysiwyg = "true";
defparam \wb_npc[29] .power_up = "low";

cyclone10lp_lcell_comb \mem_csr_data~36 (
	.dataa(\csr|io_out[29]~36_combout ),
	.datab(\csr|io_out[29]~37_combout ),
	.datac(\mem_ctrl_mem_wr~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~36_combout ),
	.cout());
defparam \mem_csr_data~36 .lut_mask = 16'hE0E0;
defparam \mem_csr_data~36 .sum_lutc_input = "datac";

dffeas \mem_csr_data[29] (
	.clk(clk_clk),
	.d(\mem_csr_data~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[29]~q ),
	.prn(vcc));
defparam \mem_csr_data[29] .is_wysiwyg = "true";
defparam \mem_csr_data[29] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[29]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~3_combout ),
	.cout());
defparam \wb_csr_data~3 .lut_mask = 16'h8888;
defparam \wb_csr_data~3 .sum_lutc_input = "datac";

dffeas \wb_csr_data[29] (
	.clk(clk_clk),
	.d(\wb_csr_data~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[29]~q ),
	.prn(vcc));
defparam \wb_csr_data[29] .is_wysiwyg = "true";
defparam \wb_csr_data[29] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[29]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~3_combout ),
	.cout());
defparam \wb_alu_out~3 .lut_mask = 16'h8888;
defparam \wb_alu_out~3 .sum_lutc_input = "datac";

dffeas \wb_alu_out[29] (
	.clk(clk_clk),
	.d(\wb_alu_out~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[29]~q ),
	.prn(vcc));
defparam \wb_alu_out[29] .is_wysiwyg = "true";
defparam \wb_alu_out[29] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[29]~9 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[29]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[29]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[29]~9_combout ),
	.cout());
defparam \_T_3543__T_3854_data[29]~9 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[29]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~37 (
	.dataa(\wb_dmem_read_data~36_combout ),
	.datab(av_readdata_pre_29),
	.datac(\wb_dmem_read_data~23_combout ),
	.datad(\wb_dmem_read_data[22]~32_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~37_combout ),
	.cout());
defparam \wb_dmem_read_data~37 .lut_mask = 16'h00AE;
defparam \wb_dmem_read_data~37 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[29] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[29]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[29] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[29] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[29]~10 (
	.dataa(\wb_npc[29]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[29]~9_combout ),
	.datad(\wb_dmem_read_data[29]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[29]~10_combout ),
	.cout());
defparam \_T_3543__T_3854_data[29]~10 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[29]~10 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a3 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[29]~10_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a3_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_a_first_bit_number = 3;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_b_first_bit_number = 3;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a3 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~5 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a3~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~5_combout ),
	.cout());
defparam \ex_rs_0~5 .lut_mask = 16'h0080;
defparam \ex_rs_0~5 .sum_lutc_input = "datac";

dffeas \ex_rs_0[29] (
	.clk(clk_clk),
	.d(\ex_rs_0~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[29]~q ),
	.prn(vcc));
defparam \ex_rs_0[29] .is_wysiwyg = "true";
defparam \ex_rs_0[29] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[29]~22 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(\ex_rs_0[29]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\wb_alu_out[29]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[29]~22_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[29]~22 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[29]~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[29]~23 (
	.dataa(av_readdata_pre_29),
	.datab(\ex_reg_rs1_bypass[2]~7_combout ),
	.datac(\ex_reg_rs1_bypass[29]~22_combout ),
	.datad(\wb_csr_data[29]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[29]~23_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[29]~23 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[29]~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[29]~24 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[29]~23_combout ),
	.datad(\mem_csr_data[29]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[29]~24_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[29]~24 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[29]~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[29]~25 (
	.dataa(\ex_reg_rs1_bypass[29]~24_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[29]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[29]~25_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[29]~25 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[29]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[29]~91 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[29]~q ),
	.datad(\ex_reg_rs1_bypass[29]~25_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[29]~91_combout ),
	.cout());
defparam \alu_io_op1[29]~91 .lut_mask = 16'h6240;
defparam \alu_io_op1[29]~91 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a3 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[29]~10_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_a_first_bit_number = 3;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_b_first_bit_number = 3;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a3 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~4 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a3~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~4_combout ),
	.cout());
defparam \ex_rs_1~4 .lut_mask = 16'h8888;
defparam \ex_rs_1~4 .sum_lutc_input = "datac";

dffeas \ex_rs_1[29] (
	.clk(clk_clk),
	.d(\ex_rs_1~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[29]~q ),
	.prn(vcc));
defparam \ex_rs_1[29] .is_wysiwyg = "true";
defparam \ex_rs_1[29] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[29]~15 (
	.dataa(\ex_reg_rs2_bypass[7]~5_combout ),
	.datab(\ex_rs_1[29]~q ),
	.datac(\ex_reg_rs2_bypass[7]~4_combout ),
	.datad(\wb_alu_out[29]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[29]~15_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[29]~15 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[29]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[29]~16 (
	.dataa(av_readdata_pre_29),
	.datab(\ex_reg_rs2_bypass[7]~5_combout ),
	.datac(\ex_reg_rs2_bypass[29]~15_combout ),
	.datad(\wb_csr_data[29]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[29]~16_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[29]~16 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[29]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[29]~17 (
	.dataa(\mem_alu_out[29]~q ),
	.datab(\ex_reg_rs2_bypass[29]~16_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[29]~17_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[29]~17 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[29]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[29]~18 (
	.dataa(\ex_reg_rs2_bypass[29]~17_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[29]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[29]~18_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[29]~18 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[29]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~4 (
	.dataa(\ex_csr_addr[9]~q ),
	.datab(\ex_ctrl_imm_type.011~q ),
	.datac(\ex_csr_addr[11]~q ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\mem_imm~4_combout ),
	.cout());
defparam \mem_imm~4 .lut_mask = 16'h88B8;
defparam \mem_imm~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[29]~73 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_reg_rs2_bypass[29]~18_combout ),
	.datad(\mem_imm~4_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[29]~73_combout ),
	.cout());
defparam \alu_io_op2[29]~73 .lut_mask = 16'hB380;
defparam \alu_io_op2[29]~73 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~24 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\alu|_T_123[29]~combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~150_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~24_combout ),
	.cout());
defparam \mem_alu_out~24 .lut_mask = 16'hDAD0;
defparam \mem_alu_out~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~25 (
	.dataa(\alu_io_op1[29]~91_combout ),
	.datab(\alu_io_op2[29]~73_combout ),
	.datac(\mem_alu_out~24_combout ),
	.datad(\alu|LessThan0~0_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~25_combout ),
	.cout());
defparam \mem_alu_out~25 .lut_mask = 16'hF08E;
defparam \mem_alu_out~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~26 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[29]~73_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~25_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~26_combout ),
	.cout());
defparam \mem_alu_out~26 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~27 (
	.dataa(\alu_io_op1[29]~91_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~26_combout ),
	.datad(\alu|ShiftRight0~130_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~27_combout ),
	.cout());
defparam \mem_alu_out~27 .lut_mask = 16'hF838;
defparam \mem_alu_out~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~28 (
	.dataa(\mem_alu_out~27_combout ),
	.datab(\alu|_T_3[29]~58_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~28_combout ),
	.cout());
defparam \mem_alu_out~28 .lut_mask = 16'h00AC;
defparam \mem_alu_out~28 .sum_lutc_input = "datac";

dffeas \mem_alu_out[29] (
	.clk(clk_clk),
	.d(\mem_alu_out~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[29]~q ),
	.prn(vcc));
defparam \mem_alu_out[29] .is_wysiwyg = "true";
defparam \mem_alu_out[29] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~27 (
	.dataa(\ex_pc[29]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~27_combout ),
	.cout());
defparam \mem_pc~27 .lut_mask = 16'h8888;
defparam \mem_pc~27 .sum_lutc_input = "datac";

dffeas \mem_pc[29] (
	.clk(clk_clk),
	.d(\mem_pc~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[29]~q ),
	.prn(vcc));
defparam \mem_pc[29] .is_wysiwyg = "true";
defparam \mem_pc[29] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~44 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\mem_imm~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_imm~44_combout ),
	.cout());
defparam \mem_imm~44 .lut_mask = 16'h8888;
defparam \mem_imm~44 .sum_lutc_input = "datac";

dffeas \mem_imm[29] (
	.clk(clk_clk),
	.d(\mem_imm~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[29]~q ),
	.prn(vcc));
defparam \mem_imm[29] .is_wysiwyg = "true";
defparam \mem_imm[29] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[29]~58 (
	.dataa(\mem_pc[29]~q ),
	.datab(\mem_imm[29]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[28]~57 ),
	.combout(\_T_3862[29]~58_combout ),
	.cout(\_T_3862[29]~59 ));
defparam \_T_3862[29]~58 .lut_mask = 16'h9617;
defparam \_T_3862[29]~58 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~91 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[29]~58_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[29]~54_combout ),
	.cin(gnd),
	.combout(\pc_cntr~91_combout ),
	.cout());
defparam \pc_cntr~91 .lut_mask = 16'h5E0E;
defparam \pc_cntr~91 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~92 (
	.dataa(\mem_alu_out[29]~q ),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~91_combout ),
	.datad(\csr|mepc[29]~q ),
	.cin(gnd),
	.combout(\pc_cntr~92_combout ),
	.cout());
defparam \pc_cntr~92 .lut_mask = 16'hF838;
defparam \pc_cntr~92 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~93 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~92_combout ),
	.datac(\csr|mtvec[29]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~93_combout ),
	.cout());
defparam \pc_cntr~93 .lut_mask = 16'h88A0;
defparam \pc_cntr~93 .sum_lutc_input = "datac";

dffeas \pc_cntr[29] (
	.clk(clk_clk),
	.d(\pc_cntr~93_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[29]~q ),
	.prn(vcc));
defparam \pc_cntr[29] .is_wysiwyg = "true";
defparam \pc_cntr[29] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~28 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[29]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~28_combout ),
	.cout());
defparam \id_pc~28 .lut_mask = 16'h8080;
defparam \id_pc~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~28 (
	.dataa(id_pc_30),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~28_combout ),
	.cout());
defparam \ex_pc~28 .lut_mask = 16'h8080;
defparam \ex_pc~28 .sum_lutc_input = "datac";

dffeas \ex_pc[30] (
	.clk(clk_clk),
	.d(\ex_pc~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[30]~q ),
	.prn(vcc));
defparam \ex_pc[30] .is_wysiwyg = "true";
defparam \ex_pc[30] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~28 (
	.dataa(\ex_pc[30]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~28_combout ),
	.cout());
defparam \mem_pc~28 .lut_mask = 16'h8888;
defparam \mem_pc~28 .sum_lutc_input = "datac";

dffeas \mem_pc[30] (
	.clk(clk_clk),
	.d(\mem_pc~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[30]~q ),
	.prn(vcc));
defparam \mem_pc[30] .is_wysiwyg = "true";
defparam \mem_pc[30] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~6 (
	.dataa(\ex_csr_addr[10]~q ),
	.datab(\ex_ctrl_imm_type.011~q ),
	.datac(\ex_csr_addr[11]~q ),
	.datad(\ex_ctrl_imm_type.101~q ),
	.cin(gnd),
	.combout(\mem_imm~6_combout ),
	.cout());
defparam \mem_imm~6 .lut_mask = 16'h88B8;
defparam \mem_imm~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_imm~45 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\mem_imm~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_imm~45_combout ),
	.cout());
defparam \mem_imm~45 .lut_mask = 16'h8888;
defparam \mem_imm~45 .sum_lutc_input = "datac";

dffeas \mem_imm[30] (
	.clk(clk_clk),
	.d(\mem_imm~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[30]~q ),
	.prn(vcc));
defparam \mem_imm[30] .is_wysiwyg = "true";
defparam \mem_imm[30] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[30]~60 (
	.dataa(\mem_pc[30]~q ),
	.datab(\mem_imm[30]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3862[29]~59 ),
	.combout(\_T_3862[30]~60_combout ),
	.cout(\_T_3862[30]~61 ));
defparam \_T_3862[30]~60 .lut_mask = 16'h698E;
defparam \_T_3862[30]~60 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \mem_csr_data~11 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[30]~45_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~11_combout ),
	.cout());
defparam \mem_csr_data~11 .lut_mask = 16'h8888;
defparam \mem_csr_data~11 .sum_lutc_input = "datac";

dffeas \mem_csr_data[30] (
	.clk(clk_clk),
	.d(\mem_csr_data~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[30]~q ),
	.prn(vcc));
defparam \mem_csr_data[30] .is_wysiwyg = "true";
defparam \mem_csr_data[30] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~4 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[30]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~4_combout ),
	.cout());
defparam \wb_csr_data~4 .lut_mask = 16'h8888;
defparam \wb_csr_data~4 .sum_lutc_input = "datac";

dffeas \wb_csr_data[30] (
	.clk(clk_clk),
	.d(\wb_csr_data~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[30]~q ),
	.prn(vcc));
defparam \wb_csr_data[30] .is_wysiwyg = "true";
defparam \wb_csr_data[30] .power_up = "low";

cyclone10lp_lcell_comb \npc[30]~56 (
	.dataa(\pc_cntr[30]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[29]~55 ),
	.combout(\npc[30]~56_combout ),
	.cout(\npc[30]~57 ));
defparam \npc[30]~56 .lut_mask = 16'hA50A;
defparam \npc[30]~56 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~4 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[30]~56_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~4_combout ),
	.cout());
defparam \id_npc~4 .lut_mask = 16'h8080;
defparam \id_npc~4 .sum_lutc_input = "datac";

dffeas \id_npc[30] (
	.clk(clk_clk),
	.d(\id_npc~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[30]~q ),
	.prn(vcc));
defparam \id_npc[30] .is_wysiwyg = "true";
defparam \id_npc[30] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~4 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[30]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~4_combout ),
	.cout());
defparam \ex_npc~4 .lut_mask = 16'h8080;
defparam \ex_npc~4 .sum_lutc_input = "datac";

dffeas \ex_npc[30] (
	.clk(clk_clk),
	.d(\ex_npc~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[30]~q ),
	.prn(vcc));
defparam \ex_npc[30] .is_wysiwyg = "true";
defparam \ex_npc[30] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~2 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[30]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~2_combout ),
	.cout());
defparam \mem_npc~2 .lut_mask = 16'h8888;
defparam \mem_npc~2 .sum_lutc_input = "datac";

dffeas \mem_npc[30] (
	.clk(clk_clk),
	.d(\mem_npc~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[30]~q ),
	.prn(vcc));
defparam \mem_npc[30] .is_wysiwyg = "true";
defparam \mem_npc[30] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[30]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~2_combout ),
	.cout());
defparam \wb_npc~2 .lut_mask = 16'h8888;
defparam \wb_npc~2 .sum_lutc_input = "datac";

dffeas \wb_npc[30] (
	.clk(clk_clk),
	.d(\wb_npc~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[30]~q ),
	.prn(vcc));
defparam \wb_npc[30] .is_wysiwyg = "true";
defparam \wb_npc[30] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~4 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[30]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~4_combout ),
	.cout());
defparam \wb_alu_out~4 .lut_mask = 16'h8888;
defparam \wb_alu_out~4 .sum_lutc_input = "datac";

dffeas \wb_alu_out[30] (
	.clk(clk_clk),
	.d(\wb_alu_out~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[30]~q ),
	.prn(vcc));
defparam \wb_alu_out[30] .is_wysiwyg = "true";
defparam \wb_alu_out[30] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[30]~11 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[30]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[30]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[30]~11_combout ),
	.cout());
defparam \_T_3543__T_3854_data[30]~11 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[30]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~38 (
	.dataa(\wb_dmem_read_data~30_combout ),
	.datab(av_readdata_pre_30),
	.datac(\wb_dmem_read_data~23_combout ),
	.datad(\wb_dmem_read_data[22]~32_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~38_combout ),
	.cout());
defparam \wb_dmem_read_data~38 .lut_mask = 16'h00AE;
defparam \wb_dmem_read_data~38 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[30] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[30]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[30] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[30] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[30]~12 (
	.dataa(\wb_csr_data[30]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[30]~11_combout ),
	.datad(\wb_dmem_read_data[30]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[30]~12_combout ),
	.cout());
defparam \_T_3543__T_3854_data[30]~12 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[30]~12 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a2 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[30]~12_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_a_first_bit_number = 2;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_b_first_bit_number = 2;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a2 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~6 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a2~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~6_combout ),
	.cout());
defparam \ex_rs_1~6 .lut_mask = 16'h8888;
defparam \ex_rs_1~6 .sum_lutc_input = "datac";

dffeas \ex_rs_1[30] (
	.clk(clk_clk),
	.d(\ex_rs_1~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[30]~q ),
	.prn(vcc));
defparam \ex_rs_1[30] .is_wysiwyg = "true";
defparam \ex_rs_1[30] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[30]~23 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_30),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[30]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[30]~23_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[30]~23 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[30]~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[30]~24 (
	.dataa(\ex_rs_1[30]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[30]~23_combout ),
	.datad(\wb_csr_data[30]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[30]~24_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[30]~24 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[30]~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[30]~25 (
	.dataa(\mem_alu_out[30]~q ),
	.datab(\ex_reg_rs2_bypass[30]~24_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[30]~25_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[30]~25 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[30]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[30]~26 (
	.dataa(\ex_reg_rs2_bypass[30]~25_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[30]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[30]~26_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[30]~26 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[30]~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[30]~75 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_reg_rs2_bypass[30]~26_combout ),
	.datad(\mem_imm~6_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[30]~75_combout ),
	.cout());
defparam \alu_io_op2[30]~75 .lut_mask = 16'hB380;
defparam \alu_io_op2[30]~75 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a2 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[30]~12_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a2_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_a_first_bit_number = 2;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_b_first_bit_number = 2;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a2 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~6 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a2~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~6_combout ),
	.cout());
defparam \ex_rs_0~6 .lut_mask = 16'h0080;
defparam \ex_rs_0~6 .sum_lutc_input = "datac";

dffeas \ex_rs_0[30] (
	.clk(clk_clk),
	.d(\ex_rs_0~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[30]~q ),
	.prn(vcc));
defparam \ex_rs_0[30] .is_wysiwyg = "true";
defparam \ex_rs_0[30] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[30]~26 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(av_readdata_pre_30),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\wb_alu_out[30]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[30]~26_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[30]~26 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[30]~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[30]~27 (
	.dataa(\ex_rs_0[30]~q ),
	.datab(\ex_reg_rs1_bypass[2]~138_combout ),
	.datac(\ex_reg_rs1_bypass[30]~26_combout ),
	.datad(\wb_csr_data[30]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[30]~27_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[30]~27 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[30]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[30]~28 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[30]~27_combout ),
	.datad(\mem_csr_data[30]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[30]~28_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[30]~28 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[30]~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[30]~29 (
	.dataa(\ex_reg_rs1_bypass[30]~28_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[30]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[30]~29_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[30]~29 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[30]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[30]~92 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[30]~q ),
	.datad(\ex_reg_rs1_bypass[30]~29_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[30]~92_combout ),
	.cout());
defparam \alu_io_op1[30]~92 .lut_mask = 16'h6240;
defparam \alu_io_op1[30]~92 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~157 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\alu_io_op2[30]~75_combout ),
	.datad(\alu_io_op1[30]~92_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~157_combout ),
	.cout());
defparam \mem_alu_out~157 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~157 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~158 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~157_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~94_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~158_combout ),
	.cout());
defparam \mem_alu_out~158 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~158 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~29 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[30]~92_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~158_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~29_combout ),
	.cout());
defparam \mem_alu_out~29 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~30 (
	.dataa(\alu_io_op2[30]~75_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~29_combout ),
	.datad(\alu|ShiftRight0~38_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~30_combout ),
	.cout());
defparam \mem_alu_out~30 .lut_mask = 16'hF838;
defparam \mem_alu_out~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~31 (
	.dataa(\mem_alu_out~30_combout ),
	.datab(\alu|_T_3[30]~60_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~31_combout ),
	.cout());
defparam \mem_alu_out~31 .lut_mask = 16'h00AC;
defparam \mem_alu_out~31 .sum_lutc_input = "datac";

dffeas \mem_alu_out[30] (
	.clk(clk_clk),
	.d(\mem_alu_out~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[30]~q ),
	.prn(vcc));
defparam \mem_alu_out[30] .is_wysiwyg = "true";
defparam \mem_alu_out[30] .power_up = "low";

cyclone10lp_lcell_comb \pc_cntr~94 (
	.dataa(\pc_cntr[19]~7_combout ),
	.datab(\mem_alu_out[30]~q ),
	.datac(\pc_cntr[19]~8_combout ),
	.datad(\npc[30]~56_combout ),
	.cin(gnd),
	.combout(\pc_cntr~94_combout ),
	.cout());
defparam \pc_cntr~94 .lut_mask = 16'hDAD0;
defparam \pc_cntr~94 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~95 (
	.dataa(\_T_3862[30]~60_combout ),
	.datab(\pc_cntr[19]~7_combout ),
	.datac(\pc_cntr~94_combout ),
	.datad(\csr|mepc[30]~q ),
	.cin(gnd),
	.combout(\pc_cntr~95_combout ),
	.cout());
defparam \pc_cntr~95 .lut_mask = 16'hF2C2;
defparam \pc_cntr~95 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~96 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~95_combout ),
	.datac(\csr|mtvec[30]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~96_combout ),
	.cout());
defparam \pc_cntr~96 .lut_mask = 16'h88A0;
defparam \pc_cntr~96 .sum_lutc_input = "datac";

dffeas \pc_cntr[30] (
	.clk(clk_clk),
	.d(\pc_cntr~96_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[30]~q ),
	.prn(vcc));
defparam \pc_cntr[30] .is_wysiwyg = "true";
defparam \pc_cntr[30] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~29 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[30]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~29_combout ),
	.cout());
defparam \id_pc~29 .lut_mask = 16'h8080;
defparam \id_pc~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_pc~29 (
	.dataa(id_pc_31),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_pc~29_combout ),
	.cout());
defparam \ex_pc~29 .lut_mask = 16'h8080;
defparam \ex_pc~29 .sum_lutc_input = "datac";

dffeas \ex_pc[31] (
	.clk(clk_clk),
	.d(\ex_pc~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_pc[31]~q ),
	.prn(vcc));
defparam \ex_pc[31] .is_wysiwyg = "true";
defparam \ex_pc[31] .power_up = "low";

cyclone10lp_lcell_comb \npc[31]~58 (
	.dataa(\pc_cntr[31]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\npc[30]~57 ),
	.combout(\npc[31]~58_combout ),
	.cout());
defparam \npc[31]~58 .lut_mask = 16'h5A5A;
defparam \npc[31]~58 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \id_npc~5 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[31]~58_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~5_combout ),
	.cout());
defparam \id_npc~5 .lut_mask = 16'h8080;
defparam \id_npc~5 .sum_lutc_input = "datac";

dffeas \id_npc[31] (
	.clk(clk_clk),
	.d(\id_npc~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[31]~q ),
	.prn(vcc));
defparam \id_npc[31] .is_wysiwyg = "true";
defparam \id_npc[31] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~5 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[31]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~5_combout ),
	.cout());
defparam \ex_npc~5 .lut_mask = 16'h8080;
defparam \ex_npc~5 .sum_lutc_input = "datac";

dffeas \ex_npc[31] (
	.clk(clk_clk),
	.d(\ex_npc~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[31]~q ),
	.prn(vcc));
defparam \ex_npc[31] .is_wysiwyg = "true";
defparam \ex_npc[31] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~3 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[31]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~3_combout ),
	.cout());
defparam \mem_npc~3 .lut_mask = 16'h8888;
defparam \mem_npc~3 .sum_lutc_input = "datac";

dffeas \mem_npc[31] (
	.clk(clk_clk),
	.d(\mem_npc~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[31]~q ),
	.prn(vcc));
defparam \mem_npc[31] .is_wysiwyg = "true";
defparam \mem_npc[31] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[31]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~3_combout ),
	.cout());
defparam \wb_npc~3 .lut_mask = 16'h8888;
defparam \wb_npc~3 .sum_lutc_input = "datac";

dffeas \wb_npc[31] (
	.clk(clk_clk),
	.d(\wb_npc~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[31]~q ),
	.prn(vcc));
defparam \wb_npc[31] .is_wysiwyg = "true";
defparam \wb_npc[31] .power_up = "low";

cyclone10lp_lcell_comb \mem_csr_data~12 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[31]~52_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~12_combout ),
	.cout());
defparam \mem_csr_data~12 .lut_mask = 16'h8888;
defparam \mem_csr_data~12 .sum_lutc_input = "datac";

dffeas \mem_csr_data[31] (
	.clk(clk_clk),
	.d(\mem_csr_data~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[31]~q ),
	.prn(vcc));
defparam \mem_csr_data[31] .is_wysiwyg = "true";
defparam \mem_csr_data[31] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~5 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[31]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~5_combout ),
	.cout());
defparam \wb_csr_data~5 .lut_mask = 16'h8888;
defparam \wb_csr_data~5 .sum_lutc_input = "datac";

dffeas \wb_csr_data[31] (
	.clk(clk_clk),
	.d(\wb_csr_data~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[31]~q ),
	.prn(vcc));
defparam \wb_csr_data[31] .is_wysiwyg = "true";
defparam \wb_csr_data[31] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~5 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_alu_out[31]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~5_combout ),
	.cout());
defparam \wb_alu_out~5 .lut_mask = 16'h8888;
defparam \wb_alu_out~5 .sum_lutc_input = "datac";

dffeas \wb_alu_out[31] (
	.clk(clk_clk),
	.d(\wb_alu_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[31]~q ),
	.prn(vcc));
defparam \wb_alu_out[31] .is_wysiwyg = "true";
defparam \wb_alu_out[31] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[31]~13 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[31]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[31]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[31]~13_combout ),
	.cout());
defparam \_T_3543__T_3854_data[31]~13 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[31]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~40 (
	.dataa(\wb_dmem_read_data~39_combout ),
	.datab(av_readdata_pre_15),
	.datac(\wb_dmem_read_data[22]~24_combout ),
	.datad(mem_alu_out_1),
	.cin(gnd),
	.combout(\wb_dmem_read_data~40_combout ),
	.cout());
defparam \wb_dmem_read_data~40 .lut_mask = 16'hAAEA;
defparam \wb_dmem_read_data~40 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~41 (
	.dataa(mem_alu_out_1),
	.datab(Equal73),
	.datac(mem_alu_out_0),
	.datad(\wb_dmem_read_data~23_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~41_combout ),
	.cout());
defparam \wb_dmem_read_data~41 .lut_mask = 16'h08FF;
defparam \wb_dmem_read_data~41 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data~42 (
	.dataa(av_readdata_pre_31),
	.datab(mem_ctrl_mem_wr01),
	.datac(\wb_dmem_read_data~40_combout ),
	.datad(\wb_dmem_read_data~41_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data~42_combout ),
	.cout());
defparam \wb_dmem_read_data~42 .lut_mask = 16'hEAC0;
defparam \wb_dmem_read_data~42 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[31] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_dmem_read_data[31]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[31] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[31] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[31]~14 (
	.dataa(\wb_npc[31]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[31]~13_combout ),
	.datad(\wb_dmem_read_data[31]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[31]~14_combout ),
	.cout());
defparam \_T_3543__T_3854_data[31]~14 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[31]~14 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a1 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[31]~14_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a1_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_a_first_bit_number = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_b_first_bit_number = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a1 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~7 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a1~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~7_combout ),
	.cout());
defparam \ex_rs_0~7 .lut_mask = 16'h0080;
defparam \ex_rs_0~7 .sum_lutc_input = "datac";

dffeas \ex_rs_0[31] (
	.clk(clk_clk),
	.d(\ex_rs_0~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[31]~q ),
	.prn(vcc));
defparam \ex_rs_0[31] .is_wysiwyg = "true";
defparam \ex_rs_0[31] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[31]~30 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(\ex_rs_0[31]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\wb_alu_out[31]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[31]~30_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[31]~30 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[31]~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[31]~31 (
	.dataa(av_readdata_pre_31),
	.datab(\ex_reg_rs1_bypass[2]~7_combout ),
	.datac(\ex_reg_rs1_bypass[31]~30_combout ),
	.datad(\wb_csr_data[31]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[31]~31_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[31]~31 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[31]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[31]~32 (
	.dataa(\_T_3634~2_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[31]~31_combout ),
	.datad(\mem_csr_data[31]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[31]~32_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[31]~32 .lut_mask = 16'hEAC0;
defparam \ex_reg_rs1_bypass[31]~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[31]~33 (
	.dataa(\ex_reg_rs1_bypass[31]~32_combout ),
	.datab(\ex_reg_rs1_bypass[0]~20_combout ),
	.datac(\mem_alu_out[31]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[31]~33_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[31]~33 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs1_bypass[31]~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[31]~93 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[31]~q ),
	.datad(\ex_reg_rs1_bypass[31]~33_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[31]~93_combout ),
	.cout());
defparam \alu_io_op1[31]~93 .lut_mask = 16'h6240;
defparam \alu_io_op1[31]~93 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a1 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[31]~14_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_a_first_bit_number = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_b_first_bit_number = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a1 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~7 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a1~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~7_combout ),
	.cout());
defparam \ex_rs_1~7 .lut_mask = 16'h8888;
defparam \ex_rs_1~7 .sum_lutc_input = "datac";

dffeas \ex_rs_1[31] (
	.clk(clk_clk),
	.d(\ex_rs_1~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[31]~q ),
	.prn(vcc));
defparam \ex_rs_1[31] .is_wysiwyg = "true";
defparam \ex_rs_1[31] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[31]~27 (
	.dataa(\ex_reg_rs2_bypass[7]~5_combout ),
	.datab(\ex_rs_1[31]~q ),
	.datac(\ex_reg_rs2_bypass[7]~4_combout ),
	.datad(\wb_alu_out[31]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[31]~27_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[31]~27 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[31]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[31]~28 (
	.dataa(av_readdata_pre_31),
	.datab(\ex_reg_rs2_bypass[7]~5_combout ),
	.datac(\ex_reg_rs2_bypass[31]~27_combout ),
	.datad(\wb_csr_data[31]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[31]~28_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[31]~28 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[31]~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[31]~29 (
	.dataa(\mem_alu_out[31]~q ),
	.datab(\ex_reg_rs2_bypass[31]~28_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[31]~29_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[31]~29 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[31]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[31]~30 (
	.dataa(\ex_reg_rs2_bypass[31]~29_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[31]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[31]~30_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[31]~30 .lut_mask = 16'hEAEA;
defparam \ex_reg_rs2_bypass[31]~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[31]~76 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_reg_rs2_bypass[31]~30_combout ),
	.datad(\mem_imm~7_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[31]~76_combout ),
	.cout());
defparam \alu_io_op2[31]~76 .lut_mask = 16'hB380;
defparam \alu_io_op2[31]~76 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~32 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\alu|_T_123[31]~combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~126_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~32_combout ),
	.cout());
defparam \mem_alu_out~32 .lut_mask = 16'hDAD0;
defparam \mem_alu_out~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~33 (
	.dataa(\alu_io_op1[31]~93_combout ),
	.datab(\alu_io_op2[31]~76_combout ),
	.datac(\mem_alu_out~32_combout ),
	.datad(\alu|LessThan0~0_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~33_combout ),
	.cout());
defparam \mem_alu_out~33 .lut_mask = 16'hF08E;
defparam \mem_alu_out~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~34 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[31]~76_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~33_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~34_combout ),
	.cout());
defparam \mem_alu_out~34 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~35 (
	.dataa(\alu_io_op1[31]~93_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~34_combout ),
	.datad(\alu|ShiftRight0~128_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~35_combout ),
	.cout());
defparam \mem_alu_out~35 .lut_mask = 16'hF838;
defparam \mem_alu_out~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~36 (
	.dataa(\mem_alu_out~35_combout ),
	.datab(\alu|_T_3[31]~62_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~36_combout ),
	.cout());
defparam \mem_alu_out~36 .lut_mask = 16'h00AC;
defparam \mem_alu_out~36 .sum_lutc_input = "datac";

dffeas \mem_alu_out[31] (
	.clk(clk_clk),
	.d(\mem_alu_out~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_alu_out[31]~q ),
	.prn(vcc));
defparam \mem_alu_out[31] .is_wysiwyg = "true";
defparam \mem_alu_out[31] .power_up = "low";

cyclone10lp_lcell_comb \mem_pc~29 (
	.dataa(\ex_pc[31]~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_pc~29_combout ),
	.cout());
defparam \mem_pc~29 .lut_mask = 16'h8888;
defparam \mem_pc~29 .sum_lutc_input = "datac";

dffeas \mem_pc[31] (
	.clk(clk_clk),
	.d(\mem_pc~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_pc[31]~q ),
	.prn(vcc));
defparam \mem_pc[31] .is_wysiwyg = "true";
defparam \mem_pc[31] .power_up = "low";

cyclone10lp_lcell_comb \mem_imm~47 (
	.dataa(\ex_csr_addr[11]~q ),
	.datab(\ex_ctrl_imm_type.101~q ),
	.datac(\mem_ctrl_mem_wr~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_imm~47_combout ),
	.cout());
defparam \mem_imm~47 .lut_mask = 16'h2020;
defparam \mem_imm~47 .sum_lutc_input = "datac";

dffeas \mem_imm[31] (
	.clk(clk_clk),
	.d(\mem_imm~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_imm[31]~q ),
	.prn(vcc));
defparam \mem_imm[31] .is_wysiwyg = "true";
defparam \mem_imm[31] .power_up = "low";

cyclone10lp_lcell_comb \_T_3862[31]~62 (
	.dataa(\mem_pc[31]~q ),
	.datab(\mem_imm[31]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\_T_3862[30]~61 ),
	.combout(\_T_3862[31]~62_combout ),
	.cout());
defparam \_T_3862[31]~62 .lut_mask = 16'h9696;
defparam \_T_3862[31]~62 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \pc_cntr~97 (
	.dataa(\pc_cntr[19]~8_combout ),
	.datab(\_T_3862[31]~62_combout ),
	.datac(\pc_cntr[19]~7_combout ),
	.datad(\npc[31]~58_combout ),
	.cin(gnd),
	.combout(\pc_cntr~97_combout ),
	.cout());
defparam \pc_cntr~97 .lut_mask = 16'h5E0E;
defparam \pc_cntr~97 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~98 (
	.dataa(\mem_alu_out[31]~q ),
	.datab(\pc_cntr[19]~8_combout ),
	.datac(\pc_cntr~97_combout ),
	.datad(\csr|mepc[31]~q ),
	.cin(gnd),
	.combout(\pc_cntr~98_combout ),
	.cout());
defparam \pc_cntr~98 .lut_mask = 16'hF838;
defparam \pc_cntr~98 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pc_cntr~99 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\pc_cntr~98_combout ),
	.datac(\csr|mtvec[31]~q ),
	.datad(\csr|io_expt~combout ),
	.cin(gnd),
	.combout(\pc_cntr~99_combout ),
	.cout());
defparam \pc_cntr~99 .lut_mask = 16'h88A0;
defparam \pc_cntr~99 .sum_lutc_input = "datac";

dffeas \pc_cntr[31] (
	.clk(clk_clk),
	.d(\pc_cntr~99_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_cntr[19]~12_combout ),
	.q(\pc_cntr[31]~q ),
	.prn(vcc));
defparam \pc_cntr[31] .is_wysiwyg = "true";
defparam \pc_cntr[31] .power_up = "low";

cyclone10lp_lcell_comb \id_pc~30 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\pc_cntr[31]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_pc~30_combout ),
	.cout());
defparam \id_pc~30 .lut_mask = 16'h8080;
defparam \id_pc~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_csr_data~8 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[1]~16_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~8_combout ),
	.cout());
defparam \mem_csr_data~8 .lut_mask = 16'h8888;
defparam \mem_csr_data~8 .sum_lutc_input = "datac";

dffeas \mem_csr_data[1] (
	.clk(clk_clk),
	.d(\mem_csr_data~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[1]~q ),
	.prn(vcc));
defparam \mem_csr_data[1] .is_wysiwyg = "true";
defparam \mem_csr_data[1] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[1]~126 (
	.dataa(\_T_3681~0_combout ),
	.datab(\_T_3681~1_combout ),
	.datac(\Equal63~0_combout ),
	.datad(\Equal62~1_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[1]~126_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[1]~126 .lut_mask = 16'h0008;
defparam \ex_reg_rs2_bypass[1]~126 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_alu_out~0 (
	.dataa(mem_alu_out_1),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~0_combout ),
	.cout());
defparam \wb_alu_out~0 .lut_mask = 16'h8888;
defparam \wb_alu_out~0 .sum_lutc_input = "datac";

dffeas \wb_alu_out[1] (
	.clk(clk_clk),
	.d(\wb_alu_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[1]~q ),
	.prn(vcc));
defparam \wb_alu_out[1] .is_wysiwyg = "true";
defparam \wb_alu_out[1] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~0 (
	.dataa(\mem_csr_data[1]~q ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~0_combout ),
	.cout());
defparam \wb_csr_data~0 .lut_mask = 16'h8888;
defparam \wb_csr_data~0 .sum_lutc_input = "datac";

dffeas \wb_csr_data[1] (
	.clk(clk_clk),
	.d(\wb_csr_data~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[1]~q ),
	.prn(vcc));
defparam \wb_csr_data[1] .is_wysiwyg = "true";
defparam \wb_csr_data[1] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[23]~0 (
	.dataa(\wb_ctrl_wb_sel.00~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\wb_ctrl_wb_sel.11~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[23]~0_combout ),
	.cout());
defparam \_T_3543__T_3854_data[23]~0 .lut_mask = 16'h00AA;
defparam \_T_3543__T_3854_data[23]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[1]~7 (
	.dataa(\wb_dmem_read_data~16_combout ),
	.datab(av_readdata_pre_17),
	.datac(gnd),
	.datad(\wb_dmem_read_data[7]~17_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data[1]~7_combout ),
	.cout());
defparam \wb_dmem_read_data[1]~7 .lut_mask = 16'hCCAA;
defparam \wb_dmem_read_data[1]~7 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[1] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data[1]~7_combout ),
	.asdata(av_readdata_pre_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\wb_dmem_read_data[7]~19_combout ),
	.sload(\wb_dmem_read_data[7]~21_combout ),
	.ena(vcc),
	.q(\wb_dmem_read_data[1]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[1] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[1] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[1]~3 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[1]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[1]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[1]~3_combout ),
	.cout());
defparam \_T_3543__T_3854_data[1]~3 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[1]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[1]~4 (
	.dataa(\_T_3543__T_3854_data[23]~0_combout ),
	.datab(\wb_ctrl_wb_sel.10~q ),
	.datac(\wb_dmem_read_data[1]~q ),
	.datad(\_T_3543__T_3854_data[1]~3_combout ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[1]~4_combout ),
	.cout());
defparam \_T_3543__T_3854_data[1]~4 .lut_mask = 16'hF100;
defparam \_T_3543__T_3854_data[1]~4 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a31 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[1]~4_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a31_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_a_first_bit_number = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_b_first_bit_number = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a31 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~2 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a31~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~2_combout ),
	.cout());
defparam \ex_rs_1~2 .lut_mask = 16'h8888;
defparam \ex_rs_1~2 .sum_lutc_input = "datac";

dffeas \ex_rs_1[1] (
	.clk(clk_clk),
	.d(\ex_rs_1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[1]~q ),
	.prn(vcc));
defparam \ex_rs_1[1] .is_wysiwyg = "true";
defparam \ex_rs_1[1] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[1]~6 (
	.dataa(\wb_csr_data[1]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_rs_1[1]~q ),
	.datad(\ex_reg_rs2_bypass[7]~5_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[1]~6_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[1]~6 .lut_mask = 16'hBBC0;
defparam \ex_reg_rs2_bypass[1]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[1]~7 (
	.dataa(av_readdata_pre_1),
	.datab(\wb_alu_out[1]~q ),
	.datac(\ex_reg_rs2_bypass[7]~4_combout ),
	.datad(\ex_reg_rs2_bypass[1]~6_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[1]~7_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[1]~7 .lut_mask = 16'hFA0C;
defparam \ex_reg_rs2_bypass[1]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[1]~8 (
	.dataa(mem_alu_out_1),
	.datab(\mem_ctrl_rf_wen~q ),
	.datac(\ex_reg_rs2_bypass[1]~7_combout ),
	.datad(\ex_reg_rs2_bypass[1]~126_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[1]~8_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[1]~8 .lut_mask = 16'hB8F0;
defparam \ex_reg_rs2_bypass[1]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[1]~9 (
	.dataa(\mem_csr_data[1]~q ),
	.datab(\mem_ctrl_csr_cmd.000~q ),
	.datac(\ex_reg_rs2_bypass[1]~126_combout ),
	.datad(\ex_reg_rs2_bypass[1]~8_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[1]~9_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[1]~9 .lut_mask = 16'hBF80;
defparam \ex_reg_rs2_bypass[1]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_alu_op2[1]~1 (
	.dataa(\csr_io_alu_op2[1]~0_combout ),
	.datab(\ex_reg_rs2_bypass[1]~9_combout ),
	.datac(\io_sw_r_ex_imm[1]~1_combout ),
	.datad(\ex_ctrl_alu_op2.10~q ),
	.cin(gnd),
	.combout(\csr_io_alu_op2[1]~1_combout ),
	.cout());
defparam \csr_io_alu_op2[1]~1 .lut_mask = 16'h88A0;
defparam \csr_io_alu_op2[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_3639~0 (
	.dataa(\mem_ctrl_rf_wen~q ),
	.datab(\Equal60~2_combout ),
	.datac(\Equal60~3_combout ),
	.datad(\Equal60~4_combout ),
	.cin(gnd),
	.combout(\_T_3639~0_combout ),
	.cout());
defparam \_T_3639~0 .lut_mask = 16'h0080;
defparam \_T_3639~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[1]~5 (
	.dataa(\_T_3639~0_combout ),
	.datab(mem_alu_out_1),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\mem_csr_data[1]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[1]~5_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[1]~5 .lut_mask = 16'hF808;
defparam \ex_reg_rs1_bypass[1]~5 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a31 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[1]~4_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a31_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_a_first_bit_number = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_b_first_bit_number = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a31 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~2 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a31~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~2_combout ),
	.cout());
defparam \ex_rs_0~2 .lut_mask = 16'h0080;
defparam \ex_rs_0~2 .sum_lutc_input = "datac";

dffeas \ex_rs_0[1] (
	.clk(clk_clk),
	.d(\ex_rs_0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[1]~q ),
	.prn(vcc));
defparam \ex_rs_0[1] .is_wysiwyg = "true";
defparam \ex_rs_0[1] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[1]~9 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(\ex_rs_0[1]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\wb_alu_out[1]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[1]~9_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[1]~9 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[1]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[1]~10 (
	.dataa(av_readdata_pre_1),
	.datab(\ex_reg_rs1_bypass[2]~7_combout ),
	.datac(\ex_reg_rs1_bypass[1]~9_combout ),
	.datad(\wb_csr_data[1]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[1]~10_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[1]~10 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[1]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[1]~11 (
	.dataa(\Equal59~1_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[1]~5_combout ),
	.datad(\ex_reg_rs1_bypass[1]~10_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[1]~11_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[1]~11 .lut_mask = 16'hDC50;
defparam \ex_reg_rs1_bypass[1]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_npc~1 (
	.dataa(id_npc_1),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~1_combout ),
	.cout());
defparam \ex_npc~1 .lut_mask = 16'h8080;
defparam \ex_npc~1 .sum_lutc_input = "datac";

dffeas \ex_npc[1] (
	.clk(clk_clk),
	.d(\ex_npc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[1]~q ),
	.prn(vcc));
defparam \ex_npc[1] .is_wysiwyg = "true";
defparam \ex_npc[1] .power_up = "low";

cyclone10lp_lcell_comb \csr_io_alu_op1[1]~7 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_reg_rs1_bypass[1]~11_combout ),
	.datad(\ex_npc[1]~q ),
	.cin(gnd),
	.combout(\csr_io_alu_op1[1]~7_combout ),
	.cout());
defparam \csr_io_alu_op1[1]~7 .lut_mask = 16'h6420;
defparam \csr_io_alu_op1[1]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~163 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\csr_io_alu_op2[1]~1_combout ),
	.datad(\csr_io_alu_op1[1]~7_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~163_combout ),
	.cout());
defparam \mem_alu_out~163 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~163 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~164 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~163_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~38_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~164_combout ),
	.cout());
defparam \mem_alu_out~164 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~164 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~3 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\csr_io_alu_op1[1]~7_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~164_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~3_combout ),
	.cout());
defparam \mem_alu_out~3 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~4 (
	.dataa(\csr_io_alu_op2[1]~1_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~3_combout ),
	.datad(\alu|ShiftRight0~94_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~4_combout ),
	.cout());
defparam \mem_alu_out~4 .lut_mask = 16'hF838;
defparam \mem_alu_out~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~7 (
	.dataa(\mem_alu_out~4_combout ),
	.datab(\alu|_T_3[1]~2_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~7_combout ),
	.cout());
defparam \mem_alu_out~7 .lut_mask = 16'h00AC;
defparam \mem_alu_out~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_csr_data~9 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[0]~24_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~9_combout ),
	.cout());
defparam \mem_csr_data~9 .lut_mask = 16'h8888;
defparam \mem_csr_data~9 .sum_lutc_input = "datac";

dffeas \mem_csr_data[0] (
	.clk(clk_clk),
	.d(\mem_csr_data~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[0]~q ),
	.prn(vcc));
defparam \mem_csr_data[0] .is_wysiwyg = "true";
defparam \mem_csr_data[0] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[0]~13 (
	.dataa(mem_alu_out_0),
	.datab(\_T_3639~0_combout ),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\mem_csr_data[0]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[0]~13_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[0]~13 .lut_mask = 16'hF808;
defparam \ex_reg_rs1_bypass[0]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_csr_data~1 (
	.dataa(\mem_csr_data[0]~q ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~1_combout ),
	.cout());
defparam \wb_csr_data~1 .lut_mask = 16'h8888;
defparam \wb_csr_data~1 .sum_lutc_input = "datac";

dffeas \wb_csr_data[0] (
	.clk(clk_clk),
	.d(\wb_csr_data~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[0]~q ),
	.prn(vcc));
defparam \wb_csr_data[0] .is_wysiwyg = "true";
defparam \wb_csr_data[0] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~1 (
	.dataa(mem_alu_out_0),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~1_combout ),
	.cout());
defparam \wb_alu_out~1 .lut_mask = 16'h8888;
defparam \wb_alu_out~1 .sum_lutc_input = "datac";

dffeas \wb_alu_out[0] (
	.clk(clk_clk),
	.d(\wb_alu_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[0]~q ),
	.prn(vcc));
defparam \wb_alu_out[0] .is_wysiwyg = "true";
defparam \wb_alu_out[0] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[0]~5 (
	.dataa(\wb_ctrl_wb_sel.00~q ),
	.datab(\wb_ctrl_wb_sel.11~q ),
	.datac(\wb_ctrl_wb_sel.10~q ),
	.datad(\wb_alu_out[0]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[0]~5_combout ),
	.cout());
defparam \_T_3543__T_3854_data[0]~5 .lut_mask = 16'hF1F0;
defparam \_T_3543__T_3854_data[0]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[0]~0 (
	.dataa(\wb_dmem_read_data~22_combout ),
	.datab(av_readdata_pre_16),
	.datac(gnd),
	.datad(\wb_dmem_read_data[7]~17_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data[0]~0_combout ),
	.cout());
defparam \wb_dmem_read_data[0]~0 .lut_mask = 16'hCCAA;
defparam \wb_dmem_read_data[0]~0 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[0] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data[0]~0_combout ),
	.asdata(av_readdata_pre_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\wb_dmem_read_data[7]~19_combout ),
	.sload(\wb_dmem_read_data[7]~21_combout ),
	.ena(vcc),
	.q(\wb_dmem_read_data[0]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[0] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[0] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[0]~6 (
	.dataa(\wb_csr_data[0]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[0]~5_combout ),
	.datad(\wb_dmem_read_data[0]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[0]~6_combout ),
	.cout());
defparam \_T_3543__T_3854_data[0]~6 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[0]~6 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a0 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[0]~6_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a0_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_a_first_bit_number = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_b_first_bit_number = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a0 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~3 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a0~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~3_combout ),
	.cout());
defparam \ex_rs_0~3 .lut_mask = 16'h0080;
defparam \ex_rs_0~3 .sum_lutc_input = "datac";

dffeas \ex_rs_0[0] (
	.clk(clk_clk),
	.d(\ex_rs_0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[0]~q ),
	.prn(vcc));
defparam \ex_rs_0[0] .is_wysiwyg = "true";
defparam \ex_rs_0[0] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[0]~14 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(av_readdata_pre_0),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\wb_alu_out[0]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[0]~14_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[0]~14 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[0]~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[0]~15 (
	.dataa(\ex_rs_0[0]~q ),
	.datab(\ex_reg_rs1_bypass[2]~138_combout ),
	.datac(\ex_reg_rs1_bypass[0]~14_combout ),
	.datad(\wb_csr_data[0]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[0]~15_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[0]~15 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[0]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[0]~16 (
	.dataa(\Equal59~1_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[0]~13_combout ),
	.datad(\ex_reg_rs1_bypass[0]~15_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[0]~16_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[0]~16 .lut_mask = 16'hDC50;
defparam \ex_reg_rs1_bypass[0]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_npc~0 (
	.dataa(id_npc_0),
	.datab(\_T_1778~combout ),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~0_combout ),
	.cout());
defparam \ex_npc~0 .lut_mask = 16'h8080;
defparam \ex_npc~0 .sum_lutc_input = "datac";

dffeas \ex_npc[0] (
	.clk(clk_clk),
	.d(\ex_npc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[0]~q ),
	.prn(vcc));
defparam \ex_npc[0] .is_wysiwyg = "true";
defparam \ex_npc[0] .power_up = "low";

cyclone10lp_lcell_comb \csr_io_alu_op1[0]~8 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_reg_rs1_bypass[0]~16_combout ),
	.datad(\ex_npc[0]~q ),
	.cin(gnd),
	.combout(\csr_io_alu_op1[0]~8_combout ),
	.cout());
defparam \csr_io_alu_op1[0]~8 .lut_mask = 16'h6420;
defparam \csr_io_alu_op1[0]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~8 (
	.dataa(\ex_ctrl_alu_func[0]~q ),
	.datab(\alu|_T_3[0]~0_combout ),
	.datac(\ex_ctrl_alu_func[1]~q ),
	.datad(\csr_io_alu_op1[0]~8_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~8_combout ),
	.cout());
defparam \mem_alu_out~8 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~9 (
	.dataa(\ex_ctrl_alu_func[2]~q ),
	.datab(\alu|_T_125~20_combout ),
	.datac(\mem_alu_out~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_alu_out~9_combout ),
	.cout());
defparam \mem_alu_out~9 .lut_mask = 16'hD8D8;
defparam \mem_alu_out~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_alu_op2[0]~2 (
	.dataa(\ex_inst[7]~q ),
	.datab(\io_sw_r_ex_imm[0]~2_combout ),
	.datac(\ex_ctrl_imm_type.001~q ),
	.datad(\ex_ctrl_alu_op2.10~q ),
	.cin(gnd),
	.combout(\csr_io_alu_op2[0]~2_combout ),
	.cout());
defparam \csr_io_alu_op2[0]~2 .lut_mask = 16'h00AC;
defparam \csr_io_alu_op2[0]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[3]~42 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\alu_io_op2[3]~42_combout ),
	.cout());
defparam \alu_io_op2[3]~42 .lut_mask = 16'h8888;
defparam \alu_io_op2[3]~42 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[0]~10 (
	.dataa(\mem_csr_data[0]~q ),
	.datab(\mem_ctrl_csr_cmd.000~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[0]~10_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[0]~10 .lut_mask = 16'h8888;
defparam \ex_reg_rs2_bypass[0]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[0]~11 (
	.dataa(\_T_3681~2_combout ),
	.datab(\Equal63~0_combout ),
	.datac(\Equal62~1_combout ),
	.datad(\ex_reg_rs2_bypass[0]~10_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[0]~11_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[0]~11 .lut_mask = 16'h0200;
defparam \ex_reg_rs2_bypass[0]~11 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a0 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[0]~6_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_a_first_bit_number = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_b_first_bit_number = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a0 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~3 (
	.dataa(\_T_3543_rtl_0|auto_generated|ram_block1a0~portbdataout ),
	.datab(\ex_rs_1[23]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~3_combout ),
	.cout());
defparam \ex_rs_1~3 .lut_mask = 16'h8888;
defparam \ex_rs_1~3 .sum_lutc_input = "datac";

dffeas \ex_rs_1[0] (
	.clk(clk_clk),
	.d(\ex_rs_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[0]~q ),
	.prn(vcc));
defparam \ex_rs_1[0] .is_wysiwyg = "true";
defparam \ex_rs_1[0] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[0]~12 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_0),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[0]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[0]~12_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[0]~12 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[0]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[0]~13 (
	.dataa(\ex_rs_1[0]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[0]~12_combout ),
	.datad(\wb_csr_data[0]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[0]~13_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[0]~13 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[0]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[0]~14 (
	.dataa(mem_alu_out_0),
	.datab(\ex_reg_rs2_bypass[0]~13_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[0]~14_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[0]~14 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[0]~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \csr_io_alu_op2[0]~3 (
	.dataa(\csr_io_alu_op2[0]~2_combout ),
	.datab(\alu_io_op2[3]~42_combout ),
	.datac(\ex_reg_rs2_bypass[0]~11_combout ),
	.datad(\ex_reg_rs2_bypass[0]~14_combout ),
	.cin(gnd),
	.combout(\csr_io_alu_op2[0]~3_combout ),
	.cout());
defparam \csr_io_alu_op2[0]~3 .lut_mask = 16'hEEEA;
defparam \csr_io_alu_op2[0]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~10 (
	.dataa(\csr_io_alu_op2[0]~3_combout ),
	.datab(\alu|ShiftRight0~126_combout ),
	.datac(\ex_ctrl_alu_func[2]~q ),
	.datad(\mem_alu_out~9_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~10_combout ),
	.cout());
defparam \mem_alu_out~10 .lut_mask = 16'hACAA;
defparam \mem_alu_out~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~11 (
	.dataa(\ex_ctrl_alu_func[3]~q ),
	.datab(\ex_ctrl_alu_func[0]~q ),
	.datac(\mem_alu_out~9_combout ),
	.datad(\mem_alu_out~10_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~11_combout ),
	.cout());
defparam \mem_alu_out~11 .lut_mask = 16'hA820;
defparam \mem_alu_out~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~12 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\mem_alu_out~11_combout ),
	.datac(\alu|io_out[0]~1_combout ),
	.datad(\ex_ctrl_alu_func[3]~q ),
	.cin(gnd),
	.combout(\mem_alu_out~12_combout ),
	.cout());
defparam \mem_alu_out~12 .lut_mask = 16'h88A8;
defparam \mem_alu_out~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_ctrl_mem_wr~8 (
	.dataa(\ex_ctrl_imm_type.001~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_ctrl_mem_wr~8_combout ),
	.cout());
defparam \mem_ctrl_mem_wr~8 .lut_mask = 16'h8888;
defparam \mem_ctrl_mem_wr~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~42 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_reg_rs2_bypass[0]~11_combout ),
	.datac(\ex_reg_rs2_bypass[0]~14_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_rs_1~42_combout ),
	.cout());
defparam \mem_rs_1~42 .lut_mask = 16'hA8A8;
defparam \mem_rs_1~42 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_csr_data~26 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[2]~150_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~26_combout ),
	.cout());
defparam \mem_csr_data~26 .lut_mask = 16'h8888;
defparam \mem_csr_data~26 .sum_lutc_input = "datac";

dffeas \mem_csr_data[2] (
	.clk(clk_clk),
	.d(\mem_csr_data~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[2]~q ),
	.prn(vcc));
defparam \mem_csr_data[2] .is_wysiwyg = "true";
defparam \mem_csr_data[2] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[2]~86 (
	.dataa(\_T_3639~0_combout ),
	.datab(mem_alu_out_2),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\mem_csr_data[2]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[2]~86_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[2]~86 .lut_mask = 16'hF808;
defparam \ex_reg_rs1_bypass[2]~86 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_csr_data~19 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~19_combout ),
	.cout());
defparam \wb_csr_data~19 .lut_mask = 16'h8888;
defparam \wb_csr_data~19 .sum_lutc_input = "datac";

dffeas \wb_csr_data[2] (
	.clk(clk_clk),
	.d(\wb_csr_data~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[2]~q ),
	.prn(vcc));
defparam \wb_csr_data[2] .is_wysiwyg = "true";
defparam \wb_csr_data[2] .power_up = "low";

cyclone10lp_lcell_comb \id_npc~19 (
	.dataa(\npc[2]~0_combout ),
	.datab(gnd),
	.datac(\_T_1778~combout ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\id_npc~19_combout ),
	.cout());
defparam \id_npc~19 .lut_mask = 16'hAFFF;
defparam \id_npc~19 .sum_lutc_input = "datac";

dffeas \id_npc[2] (
	.clk(clk_clk),
	.d(\id_npc~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[2]~q ),
	.prn(vcc));
defparam \id_npc[2] .is_wysiwyg = "true";
defparam \id_npc[2] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~19 (
	.dataa(\id_npc[2]~q ),
	.datab(gnd),
	.datac(\_T_1778~combout ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\ex_npc~19_combout ),
	.cout());
defparam \ex_npc~19 .lut_mask = 16'hAFFF;
defparam \ex_npc~19 .sum_lutc_input = "datac";

dffeas \ex_npc[2] (
	.clk(clk_clk),
	.d(\ex_npc~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[2]~q ),
	.prn(vcc));
defparam \ex_npc[2] .is_wysiwyg = "true";
defparam \ex_npc[2] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~17 (
	.dataa(\ex_npc[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_npc~17_combout ),
	.cout());
defparam \mem_npc~17 .lut_mask = 16'hAAFF;
defparam \mem_npc~17 .sum_lutc_input = "datac";

dffeas \mem_npc[2] (
	.clk(clk_clk),
	.d(\mem_npc~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[2]~q ),
	.prn(vcc));
defparam \mem_npc[2] .is_wysiwyg = "true";
defparam \mem_npc[2] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~17 (
	.dataa(\mem_npc[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\wb_npc~17_combout ),
	.cout());
defparam \wb_npc~17 .lut_mask = 16'hAAFF;
defparam \wb_npc~17 .sum_lutc_input = "datac";

dffeas \wb_npc[2] (
	.clk(clk_clk),
	.d(\wb_npc~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[2]~q ),
	.prn(vcc));
defparam \wb_npc[2] .is_wysiwyg = "true";
defparam \wb_npc[2] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~19 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(mem_alu_out_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~19_combout ),
	.cout());
defparam \wb_alu_out~19 .lut_mask = 16'h8888;
defparam \wb_alu_out~19 .sum_lutc_input = "datac";

dffeas \wb_alu_out[2] (
	.clk(clk_clk),
	.d(\wb_alu_out~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[2]~q ),
	.prn(vcc));
defparam \wb_alu_out[2] .is_wysiwyg = "true";
defparam \wb_alu_out[2] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[2]~41 (
	.dataa(\_T_3543__T_3854_data[23]~2_combout ),
	.datab(\wb_npc[2]~q ),
	.datac(\_T_3543__T_3854_data[23]~1_combout ),
	.datad(\wb_alu_out[2]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[2]~41_combout ),
	.cout());
defparam \_T_3543__T_3854_data[2]~41 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[2]~41 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[2]~6 (
	.dataa(\wb_dmem_read_data~52_combout ),
	.datab(av_readdata_pre_18),
	.datac(gnd),
	.datad(\wb_dmem_read_data[7]~17_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data[2]~6_combout ),
	.cout());
defparam \wb_dmem_read_data[2]~6 .lut_mask = 16'hCCAA;
defparam \wb_dmem_read_data[2]~6 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[2] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data[2]~6_combout ),
	.asdata(av_readdata_pre_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\wb_dmem_read_data[7]~19_combout ),
	.sload(\wb_dmem_read_data[7]~21_combout ),
	.ena(vcc),
	.q(\wb_dmem_read_data[2]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[2] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[2] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[2]~42 (
	.dataa(\wb_csr_data[2]~q ),
	.datab(\_T_3543__T_3854_data[23]~2_combout ),
	.datac(\_T_3543__T_3854_data[2]~41_combout ),
	.datad(\wb_dmem_read_data[2]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[2]~42_combout ),
	.cout());
defparam \_T_3543__T_3854_data[2]~42 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[2]~42 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a30 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[2]~42_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a30_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_a_first_bit_number = 30;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_b_first_bit_number = 30;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a30 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~21 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a30~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~21_combout ),
	.cout());
defparam \ex_rs_0~21 .lut_mask = 16'h0080;
defparam \ex_rs_0~21 .sum_lutc_input = "datac";

dffeas \ex_rs_0[2] (
	.clk(clk_clk),
	.d(\ex_rs_0~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[2]~q ),
	.prn(vcc));
defparam \ex_rs_0[2] .is_wysiwyg = "true";
defparam \ex_rs_0[2] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[2]~87 (
	.dataa(\ex_reg_rs1_bypass[2]~138_combout ),
	.datab(av_readdata_pre_2),
	.datac(\ex_reg_rs1_bypass[2]~7_combout ),
	.datad(\wb_alu_out[2]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[2]~87_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[2]~87 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[2]~87 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[2]~88 (
	.dataa(\ex_rs_0[2]~q ),
	.datab(\ex_reg_rs1_bypass[2]~138_combout ),
	.datac(\ex_reg_rs1_bypass[2]~87_combout ),
	.datad(\wb_csr_data[2]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[2]~88_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[2]~88 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[2]~88 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[2]~89 (
	.dataa(\Equal59~1_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[2]~86_combout ),
	.datad(\ex_reg_rs1_bypass[2]~88_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[2]~89_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[2]~89 .lut_mask = 16'hDC50;
defparam \ex_reg_rs1_bypass[2]~89 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[2]~107 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[2]~q ),
	.datad(\ex_reg_rs1_bypass[2]~89_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[2]~107_combout ),
	.cout());
defparam \alu_io_op1[2]~107 .lut_mask = 16'h6240;
defparam \alu_io_op1[2]~107 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[2]~77 (
	.dataa(\_T_3681~3_combout ),
	.datab(\mem_csr_data[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[2]~77_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[2]~77 .lut_mask = 16'h8888;
defparam \ex_reg_rs2_bypass[2]~77 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a30 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[2]~42_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a30_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_a_first_bit_number = 30;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_b_first_bit_number = 30;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a30 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~21 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a30~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~21_combout ),
	.cout());
defparam \ex_rs_1~21 .lut_mask = 16'h8888;
defparam \ex_rs_1~21 .sum_lutc_input = "datac";

dffeas \ex_rs_1[2] (
	.clk(clk_clk),
	.d(\ex_rs_1~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[2]~q ),
	.prn(vcc));
defparam \ex_rs_1[2] .is_wysiwyg = "true";
defparam \ex_rs_1[2] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[2]~78 (
	.dataa(\ex_reg_rs2_bypass[7]~4_combout ),
	.datab(av_readdata_pre_2),
	.datac(\ex_reg_rs2_bypass[7]~5_combout ),
	.datad(\wb_alu_out[2]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[2]~78_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[2]~78 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs2_bypass[2]~78 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[2]~79 (
	.dataa(\ex_rs_1[2]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_reg_rs2_bypass[2]~78_combout ),
	.datad(\wb_csr_data[2]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[2]~79_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[2]~79 .lut_mask = 16'hF838;
defparam \ex_reg_rs2_bypass[2]~79 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[2]~80 (
	.dataa(mem_alu_out_2),
	.datab(\ex_reg_rs2_bypass[2]~79_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[2]~80_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[2]~80 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[2]~80 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[2]~63 (
	.dataa(\io_sw_r_ex_imm[2]~6_combout ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_reg_rs2_bypass[2]~77_combout ),
	.datad(\ex_reg_rs2_bypass[2]~80_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[2]~63_combout ),
	.cout());
defparam \alu_io_op2[2]~63 .lut_mask = 16'hEEE2;
defparam \alu_io_op2[2]~63 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[2]~91 (
	.dataa(\ex_ctrl_alu_op2.01~q ),
	.datab(\ex_ctrl_alu_op2.10~q ),
	.datac(\ex_ctrl_imm_type.011~q ),
	.datad(\alu_io_op2[2]~63_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[2]~91_combout ),
	.cout());
defparam \alu_io_op2[2]~91 .lut_mask = 16'h8B00;
defparam \alu_io_op2[2]~91 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~13 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\alu|_T_123[2]~combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~130_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~13_combout ),
	.cout());
defparam \mem_alu_out~13 .lut_mask = 16'hDAD0;
defparam \mem_alu_out~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~14 (
	.dataa(\alu_io_op1[2]~107_combout ),
	.datab(\alu_io_op2[2]~91_combout ),
	.datac(\mem_alu_out~13_combout ),
	.datad(\alu|LessThan0~0_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~14_combout ),
	.cout());
defparam \mem_alu_out~14 .lut_mask = 16'hF08E;
defparam \mem_alu_out~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~15 (
	.dataa(\mem_alu_out[26]~1_combout ),
	.datab(\alu_io_op2[2]~91_combout ),
	.datac(\mem_alu_out[26]~0_combout ),
	.datad(\mem_alu_out~14_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~15_combout ),
	.cout());
defparam \mem_alu_out~15 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~16 (
	.dataa(\alu_io_op1[2]~107_combout ),
	.datab(\mem_alu_out[26]~1_combout ),
	.datac(\mem_alu_out~15_combout ),
	.datad(\alu|ShiftRight0~150_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~16_combout ),
	.cout());
defparam \mem_alu_out~16 .lut_mask = 16'hF838;
defparam \mem_alu_out~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~17 (
	.dataa(\mem_alu_out~16_combout ),
	.datab(\alu|_T_3[2]~4_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~17_combout ),
	.cout());
defparam \mem_alu_out~17 .lut_mask = 16'h00AC;
defparam \mem_alu_out~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_csr_data~27 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\csr|io_out[3]~159_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_csr_data~27_combout ),
	.cout());
defparam \mem_csr_data~27 .lut_mask = 16'h8888;
defparam \mem_csr_data~27 .sum_lutc_input = "datac";

dffeas \mem_csr_data[3] (
	.clk(clk_clk),
	.d(\mem_csr_data~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_csr_data[3]~q ),
	.prn(vcc));
defparam \mem_csr_data[3] .is_wysiwyg = "true";
defparam \mem_csr_data[3] .power_up = "low";

cyclone10lp_lcell_comb \wb_alu_out~20 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(mem_alu_out_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_alu_out~20_combout ),
	.cout());
defparam \wb_alu_out~20 .lut_mask = 16'h8888;
defparam \wb_alu_out~20 .sum_lutc_input = "datac";

dffeas \wb_alu_out[3] (
	.clk(clk_clk),
	.d(\wb_alu_out~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_alu_out[3]~q ),
	.prn(vcc));
defparam \wb_alu_out[3] .is_wysiwyg = "true";
defparam \wb_alu_out[3] .power_up = "low";

cyclone10lp_lcell_comb \wb_csr_data~20 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_csr_data[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_csr_data~20_combout ),
	.cout());
defparam \wb_csr_data~20 .lut_mask = 16'h8888;
defparam \wb_csr_data~20 .sum_lutc_input = "datac";

dffeas \wb_csr_data[3] (
	.clk(clk_clk),
	.d(\wb_csr_data~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_csr_data[3]~q ),
	.prn(vcc));
defparam \wb_csr_data[3] .is_wysiwyg = "true";
defparam \wb_csr_data[3] .power_up = "low";

cyclone10lp_lcell_comb \id_npc~20 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\npc[3]~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\id_npc~20_combout ),
	.cout());
defparam \id_npc~20 .lut_mask = 16'h8080;
defparam \id_npc~20 .sum_lutc_input = "datac";

dffeas \id_npc[3] (
	.clk(clk_clk),
	.d(\id_npc~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\id_pc[7]~0_combout ),
	.q(\id_npc[3]~q ),
	.prn(vcc));
defparam \id_npc[3] .is_wysiwyg = "true";
defparam \id_npc[3] .power_up = "low";

cyclone10lp_lcell_comb \ex_npc~20 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\id_npc[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_npc~20_combout ),
	.cout());
defparam \ex_npc~20 .lut_mask = 16'h8080;
defparam \ex_npc~20 .sum_lutc_input = "datac";

dffeas \ex_npc[3] (
	.clk(clk_clk),
	.d(\ex_npc~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_npc[3]~q ),
	.prn(vcc));
defparam \ex_npc[3] .is_wysiwyg = "true";
defparam \ex_npc[3] .power_up = "low";

cyclone10lp_lcell_comb \mem_npc~18 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_npc[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_npc~18_combout ),
	.cout());
defparam \mem_npc~18 .lut_mask = 16'h8888;
defparam \mem_npc~18 .sum_lutc_input = "datac";

dffeas \mem_npc[3] (
	.clk(clk_clk),
	.d(\mem_npc~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_npc[3]~q ),
	.prn(vcc));
defparam \mem_npc[3] .is_wysiwyg = "true";
defparam \mem_npc[3] .power_up = "low";

cyclone10lp_lcell_comb \wb_npc~18 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\mem_npc[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wb_npc~18_combout ),
	.cout());
defparam \wb_npc~18 .lut_mask = 16'h8888;
defparam \wb_npc~18 .sum_lutc_input = "datac";

dffeas \wb_npc[3] (
	.clk(clk_clk),
	.d(\wb_npc~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wb_npc[3]~q ),
	.prn(vcc));
defparam \wb_npc[3] .is_wysiwyg = "true";
defparam \wb_npc[3] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[3]~43 (
	.dataa(\_T_3543__T_3854_data[23]~1_combout ),
	.datab(\wb_csr_data[3]~q ),
	.datac(\_T_3543__T_3854_data[23]~2_combout ),
	.datad(\wb_alu_out[3]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[3]~43_combout ),
	.cout());
defparam \_T_3543__T_3854_data[3]~43 .lut_mask = 16'hE5E0;
defparam \_T_3543__T_3854_data[3]~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wb_dmem_read_data[3]~5 (
	.dataa(\wb_dmem_read_data~56_combout ),
	.datab(av_readdata_pre_19),
	.datac(gnd),
	.datad(\wb_dmem_read_data[7]~17_combout ),
	.cin(gnd),
	.combout(\wb_dmem_read_data[3]~5_combout ),
	.cout());
defparam \wb_dmem_read_data[3]~5 .lut_mask = 16'hCCAA;
defparam \wb_dmem_read_data[3]~5 .sum_lutc_input = "datac";

dffeas \wb_dmem_read_data[3] (
	.clk(clk_clk),
	.d(\wb_dmem_read_data[3]~5_combout ),
	.asdata(av_readdata_pre_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\wb_dmem_read_data[7]~19_combout ),
	.sload(\wb_dmem_read_data[7]~21_combout ),
	.ena(vcc),
	.q(\wb_dmem_read_data[3]~q ),
	.prn(vcc));
defparam \wb_dmem_read_data[3] .is_wysiwyg = "true";
defparam \wb_dmem_read_data[3] .power_up = "low";

cyclone10lp_lcell_comb \_T_3543__T_3854_data[3]~44 (
	.dataa(\wb_npc[3]~q ),
	.datab(\_T_3543__T_3854_data[23]~1_combout ),
	.datac(\_T_3543__T_3854_data[3]~43_combout ),
	.datad(\wb_dmem_read_data[3]~q ),
	.cin(gnd),
	.combout(\_T_3543__T_3854_data[3]~44_combout ),
	.cout());
defparam \_T_3543__T_3854_data[3]~44 .lut_mask = 16'hF838;
defparam \_T_3543__T_3854_data[3]~44 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_0|auto_generated|ram_block1a29 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[3]~44_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~20_combout ,\id_inst~16_combout ,\id_inst~18_combout ,\id_inst~12_combout ,\id_inst~14_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_0|auto_generated|ram_block1a29_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_0|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .operation_mode = "dual_port";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_a_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_a_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_a_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_a_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_a_first_bit_number = 29;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_a_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_b_address_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_b_address_width = 5;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_b_data_width = 1;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_b_first_address = 0;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_b_first_bit_number = 29;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_b_last_address = 31;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_0|auto_generated|ram_block1a29 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_1~22 (
	.dataa(\ex_rs_1[23]~1_combout ),
	.datab(\_T_3543_rtl_0|auto_generated|ram_block1a29~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ex_rs_1~22_combout ),
	.cout());
defparam \ex_rs_1~22 .lut_mask = 16'h8888;
defparam \ex_rs_1~22 .sum_lutc_input = "datac";

dffeas \ex_rs_1[3] (
	.clk(clk_clk),
	.d(\ex_rs_1~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_1[3]~q ),
	.prn(vcc));
defparam \ex_rs_1[3] .is_wysiwyg = "true";
defparam \ex_rs_1[3] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[3]~81 (
	.dataa(\wb_csr_data[3]~q ),
	.datab(\ex_reg_rs2_bypass[7]~4_combout ),
	.datac(\ex_rs_1[3]~q ),
	.datad(\ex_reg_rs2_bypass[7]~5_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[3]~81_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[3]~81 .lut_mask = 16'hBBC0;
defparam \ex_reg_rs2_bypass[3]~81 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[3]~82 (
	.dataa(av_readdata_pre_3),
	.datab(\wb_alu_out[3]~q ),
	.datac(\ex_reg_rs2_bypass[7]~4_combout ),
	.datad(\ex_reg_rs2_bypass[3]~81_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[3]~82_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[3]~82 .lut_mask = 16'hFA0C;
defparam \ex_reg_rs2_bypass[3]~82 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[3]~64 (
	.dataa(mem_alu_out_3),
	.datab(\_T_3686~0_combout ),
	.datac(\ex_reg_rs2_bypass[3]~82_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\alu_io_op2[3]~64_combout ),
	.cout());
defparam \alu_io_op2[3]~64 .lut_mask = 16'hB8B8;
defparam \alu_io_op2[3]~64 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[3]~65 (
	.dataa(\alu_io_op2[3]~42_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[3]~q ),
	.datad(\alu_io_op2[3]~64_combout ),
	.cin(gnd),
	.combout(\alu_io_op2[3]~65_combout ),
	.cout());
defparam \alu_io_op2[3]~65 .lut_mask = 16'hA280;
defparam \alu_io_op2[3]~65 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op2[3]~66 (
	.dataa(\alu_io_op2[3]~65_combout ),
	.datab(\io_sw_r_ex_imm[3]~8_combout ),
	.datac(\ex_ctrl_alu_op2.10~q ),
	.datad(\ex_ctrl_imm_type.011~q ),
	.cin(gnd),
	.combout(\alu_io_op2[3]~66_combout ),
	.cout());
defparam \alu_io_op2[3]~66 .lut_mask = 16'hAAAE;
defparam \alu_io_op2[3]~66 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[3]~94 (
	.dataa(\_T_3639~0_combout ),
	.datab(mem_alu_out_3),
	.datac(\csr_io_in[0]~0_combout ),
	.datad(\mem_csr_data[3]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[3]~94_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[3]~94 .lut_mask = 16'hF808;
defparam \ex_reg_rs1_bypass[3]~94 .sum_lutc_input = "datac";

cyclone10lp_ram_block \_T_3543_rtl_1|auto_generated|ram_block1a29 (
	.portawe(\_T_3543__T_3854_en~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(!clk_clk),
	.clk1(clk_clk),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\_T_3543__T_3854_data[3]~44_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wb_reg_waddr[4]~q ,\wb_reg_waddr[3]~q ,\wb_reg_waddr[2]~q ,\wb_reg_waddr[1]~q ,\wb_reg_waddr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\id_inst~10_combout ,\id_inst~6_combout ,\id_inst~8_combout ,\id_inst~2_combout ,\id_inst~4_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\_T_3543_rtl_1|auto_generated|ram_block1a29_PORTBDATAOUT_bus ));
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .data_interleave_offset_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .data_interleave_width_in_bits = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .logical_ram_name = "kyogenrv_fpga_avalonMM:kyogenrv_0|KyogenRVCpu:krv|altsyncram:_T_3543_rtl_1|altsyncram_dvc1:auto_generated|ALTSYNCRAM";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .mixed_port_feed_through_mode = "dont_care";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .operation_mode = "dual_port";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_a_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_a_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_a_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_a_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_a_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_a_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_a_first_bit_number = 29;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_a_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_a_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_a_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_b_address_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_b_address_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_b_address_width = 5;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_b_data_out_clear = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_b_data_out_clock = "none";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_b_data_width = 1;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_b_first_address = 0;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_b_first_bit_number = 29;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_b_last_address = 31;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_b_logical_ram_depth = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_b_logical_ram_width = 32;
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .port_b_read_enable_clock = "clock1";
defparam \_T_3543_rtl_1|auto_generated|ram_block1a29 .ram_block_type = "auto";

cyclone10lp_lcell_comb \ex_rs_0~23 (
	.dataa(\_T_1778~combout ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(\_T_3543_rtl_1|auto_generated|ram_block1a29~portbdataout ),
	.datad(\ex_rs_0[3]~1_combout ),
	.cin(gnd),
	.combout(\ex_rs_0~23_combout ),
	.cout());
defparam \ex_rs_0~23 .lut_mask = 16'h0080;
defparam \ex_rs_0~23 .sum_lutc_input = "datac";

dffeas \ex_rs_0[3] (
	.clk(clk_clk),
	.d(\ex_rs_0~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_rs_0[3]~q ),
	.prn(vcc));
defparam \ex_rs_0[3] .is_wysiwyg = "true";
defparam \ex_rs_0[3] .power_up = "low";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[3]~95 (
	.dataa(\ex_reg_rs1_bypass[2]~7_combout ),
	.datab(\ex_rs_0[3]~q ),
	.datac(\ex_reg_rs1_bypass[2]~138_combout ),
	.datad(\wb_alu_out[3]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[3]~95_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[3]~95 .lut_mask = 16'hE5E0;
defparam \ex_reg_rs1_bypass[3]~95 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[3]~96 (
	.dataa(av_readdata_pre_3),
	.datab(\ex_reg_rs1_bypass[2]~7_combout ),
	.datac(\ex_reg_rs1_bypass[3]~95_combout ),
	.datad(\wb_csr_data[3]~q ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[3]~96_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[3]~96 .lut_mask = 16'hF838;
defparam \ex_reg_rs1_bypass[3]~96 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs1_bypass[3]~97 (
	.dataa(\Equal59~1_combout ),
	.datab(\ex_reg_rs1_bypass[0]~4_combout ),
	.datac(\ex_reg_rs1_bypass[3]~94_combout ),
	.datad(\ex_reg_rs1_bypass[3]~96_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs1_bypass[3]~97_combout ),
	.cout());
defparam \ex_reg_rs1_bypass[3]~97 .lut_mask = 16'hDC50;
defparam \ex_reg_rs1_bypass[3]~97 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \alu_io_op1[3]~109 (
	.dataa(\ex_ctrl_alu_op1[0]~q ),
	.datab(\ex_ctrl_alu_op1[1]~q ),
	.datac(\ex_pc[3]~q ),
	.datad(\ex_reg_rs1_bypass[3]~97_combout ),
	.cin(gnd),
	.combout(\alu_io_op1[3]~109_combout ),
	.cout());
defparam \alu_io_op1[3]~109 .lut_mask = 16'h6240;
defparam \alu_io_op1[3]~109 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~161 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out[26]~2_combout ),
	.datac(\alu_io_op2[3]~66_combout ),
	.datad(\alu_io_op1[3]~109_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~161_combout ),
	.cout());
defparam \mem_alu_out~161 .lut_mask = 16'h7BB2;
defparam \mem_alu_out~161 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~162 (
	.dataa(\alu|LessThan0~0_combout ),
	.datab(\mem_alu_out~161_combout ),
	.datac(\mem_alu_out[26]~2_combout ),
	.datad(\alu|ShiftRight0~152_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~162_combout ),
	.cout());
defparam \mem_alu_out~162 .lut_mask = 16'hCCC4;
defparam \mem_alu_out~162 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~18 (
	.dataa(\mem_alu_out[26]~0_combout ),
	.datab(\alu_io_op1[3]~109_combout ),
	.datac(\mem_alu_out[26]~1_combout ),
	.datad(\mem_alu_out~162_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~18_combout ),
	.cout());
defparam \mem_alu_out~18 .lut_mask = 16'hE5E0;
defparam \mem_alu_out~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~19 (
	.dataa(\alu_io_op2[3]~66_combout ),
	.datab(\mem_alu_out[26]~0_combout ),
	.datac(\mem_alu_out~18_combout ),
	.datad(\alu|ShiftRight0~167_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~19_combout ),
	.cout());
defparam \mem_alu_out~19 .lut_mask = 16'hF838;
defparam \mem_alu_out~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_alu_out~20 (
	.dataa(\mem_alu_out~19_combout ),
	.datab(\alu|_T_3[3]~6_combout ),
	.datac(\mem_alu_out[26]~5_combout ),
	.datad(\mem_alu_out[26]~6_combout ),
	.cin(gnd),
	.combout(\mem_alu_out~20_combout ),
	.cout());
defparam \mem_alu_out~20 .lut_mask = 16'h00AC;
defparam \mem_alu_out~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~43 (
	.dataa(\ex_reg_rs2_bypass[1]~9_combout ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_rs_1~43_combout ),
	.cout());
defparam \mem_rs_1~43 .lut_mask = 16'h8888;
defparam \mem_rs_1~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~53 (
	.dataa(\_T_3681~3_combout ),
	.datab(\mem_csr_data[2]~q ),
	.datac(\mem_ctrl_mem_wr~7_combout ),
	.datad(\ex_reg_rs2_bypass[2]~80_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~53_combout ),
	.cout());
defparam \mem_rs_1~53 .lut_mask = 16'hF080;
defparam \mem_rs_1~53 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[3]~124 (
	.dataa(mem_alu_out_3),
	.datab(\ex_reg_rs2_bypass[3]~82_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[3]~124_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[3]~124 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[3]~124 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~44 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_reg_rs2_bypass[3]~124_combout ),
	.datac(\_T_3681~3_combout ),
	.datad(\mem_csr_data[3]~q ),
	.cin(gnd),
	.combout(\mem_rs_1~44_combout ),
	.cout());
defparam \mem_rs_1~44 .lut_mask = 16'hA888;
defparam \mem_rs_1~44 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_reg_rs2_bypass[4]~125 (
	.dataa(\mem_alu_out[4]~q ),
	.datab(\ex_reg_rs2_bypass[4]~76_combout ),
	.datac(\_T_3686~0_combout ),
	.datad(\_T_3681~3_combout ),
	.cin(gnd),
	.combout(\ex_reg_rs2_bypass[4]~125_combout ),
	.cout());
defparam \ex_reg_rs2_bypass[4]~125 .lut_mask = 16'h00AC;
defparam \ex_reg_rs2_bypass[4]~125 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~45 (
	.dataa(\mem_ctrl_mem_wr~7_combout ),
	.datab(\ex_reg_rs2_bypass[4]~125_combout ),
	.datac(\_T_3681~3_combout ),
	.datad(\mem_csr_data[4]~q ),
	.cin(gnd),
	.combout(\mem_rs_1~45_combout ),
	.cout());
defparam \mem_rs_1~45 .lut_mask = 16'hA888;
defparam \mem_rs_1~45 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~46 (
	.dataa(\ex_reg_rs2_bypass[5]~85_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[5]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~46_combout ),
	.cout());
defparam \mem_rs_1~46 .lut_mask = 16'hEA00;
defparam \mem_rs_1~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~47 (
	.dataa(\ex_reg_rs2_bypass[6]~88_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[6]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~47_combout ),
	.cout());
defparam \mem_rs_1~47 .lut_mask = 16'hEA00;
defparam \mem_rs_1~47 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~48 (
	.dataa(\ex_reg_rs2_bypass[7]~91_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[7]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~48_combout ),
	.cout());
defparam \mem_rs_1~48 .lut_mask = 16'hEA00;
defparam \mem_rs_1~48 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~49 (
	.dataa(\ex_reg_rs2_bypass[8]~36_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[8]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~49_combout ),
	.cout());
defparam \mem_rs_1~49 .lut_mask = 16'hEA00;
defparam \mem_rs_1~49 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~50 (
	.dataa(\ex_reg_rs2_bypass[9]~33_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[9]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~50_combout ),
	.cout());
defparam \mem_rs_1~50 .lut_mask = 16'hEA00;
defparam \mem_rs_1~50 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~51 (
	.dataa(\ex_reg_rs2_bypass[10]~39_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[10]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~51_combout ),
	.cout());
defparam \mem_rs_1~51 .lut_mask = 16'hEA00;
defparam \mem_rs_1~51 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~52 (
	.dataa(\ex_reg_rs2_bypass[11]~42_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[11]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~52_combout ),
	.cout());
defparam \mem_rs_1~52 .lut_mask = 16'hEA00;
defparam \mem_rs_1~52 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~54 (
	.dataa(\ex_reg_rs2_bypass[12]~49_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[12]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~54_combout ),
	.cout());
defparam \mem_rs_1~54 .lut_mask = 16'hEA00;
defparam \mem_rs_1~54 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~55 (
	.dataa(\ex_reg_rs2_bypass[13]~45_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[13]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~55_combout ),
	.cout());
defparam \mem_rs_1~55 .lut_mask = 16'hEA00;
defparam \mem_rs_1~55 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~56 (
	.dataa(\ex_reg_rs2_bypass[14]~53_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[14]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~56_combout ),
	.cout());
defparam \mem_rs_1~56 .lut_mask = 16'hEA00;
defparam \mem_rs_1~56 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~57 (
	.dataa(\ex_reg_rs2_bypass[15]~57_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[15]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~57_combout ),
	.cout());
defparam \mem_rs_1~57 .lut_mask = 16'hEA00;
defparam \mem_rs_1~57 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~58 (
	.dataa(\ex_reg_rs2_bypass[16]~65_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[16]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~58_combout ),
	.cout());
defparam \mem_rs_1~58 .lut_mask = 16'hEA00;
defparam \mem_rs_1~58 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~59 (
	.dataa(\ex_reg_rs2_bypass[17]~61_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[17]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~59_combout ),
	.cout());
defparam \mem_rs_1~59 .lut_mask = 16'hEA00;
defparam \mem_rs_1~59 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~60 (
	.dataa(\ex_reg_rs2_bypass[18]~69_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[18]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~60_combout ),
	.cout());
defparam \mem_rs_1~60 .lut_mask = 16'hEA00;
defparam \mem_rs_1~60 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~61 (
	.dataa(\ex_reg_rs2_bypass[19]~73_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[19]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~61_combout ),
	.cout());
defparam \mem_rs_1~61 .lut_mask = 16'hEA00;
defparam \mem_rs_1~61 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~62 (
	.dataa(\ex_reg_rs2_bypass[20]~98_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[20]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~62_combout ),
	.cout());
defparam \mem_rs_1~62 .lut_mask = 16'hEA00;
defparam \mem_rs_1~62 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~63 (
	.dataa(\ex_reg_rs2_bypass[21]~94_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[21]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~63_combout ),
	.cout());
defparam \mem_rs_1~63 .lut_mask = 16'hEA00;
defparam \mem_rs_1~63 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~64 (
	.dataa(\ex_reg_rs2_bypass[22]~102_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[22]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~64_combout ),
	.cout());
defparam \mem_rs_1~64 .lut_mask = 16'hEA00;
defparam \mem_rs_1~64 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~65 (
	.dataa(\ex_reg_rs2_bypass[23]~106_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[23]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~65_combout ),
	.cout());
defparam \mem_rs_1~65 .lut_mask = 16'hEA00;
defparam \mem_rs_1~65 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mem_wr~12 (
	.dataa(\ex_ctrl_mem_wr~8_combout ),
	.datab(\ex_ctrl_mask_type~0_combout ),
	.datac(\_GEN_15~2_combout ),
	.datad(\ex_ctrl_mem_wr~9_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_mem_wr~12_combout ),
	.cout());
defparam \ex_ctrl_mem_wr~12 .lut_mask = 16'hFF40;
defparam \ex_ctrl_mem_wr~12 .sum_lutc_input = "datac";

dffeas \ex_ctrl_mem_wr.00 (
	.clk(clk_clk),
	.d(\ex_ctrl_mem_wr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_mem_wr.00~q ),
	.prn(vcc));
defparam \ex_ctrl_mem_wr.00 .is_wysiwyg = "true";
defparam \ex_ctrl_mem_wr.00 .power_up = "low";

cyclone10lp_lcell_comb \mem_ctrl_mem_wr~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\mem_ctrl_mem_wr~7_combout ),
	.datad(\ex_ctrl_mem_wr.00~q ),
	.cin(gnd),
	.combout(\mem_ctrl_mem_wr~9_combout ),
	.cout());
defparam \mem_ctrl_mem_wr~9 .lut_mask = 16'hF000;
defparam \mem_ctrl_mem_wr~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \w_req~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\w_req~0_combout ),
	.cout());
defparam \w_req~0 .lut_mask = 16'h5555;
defparam \w_req~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mem_wr~11 (
	.dataa(\id_inst[14]~q ),
	.datab(\id_inst[12]~q ),
	.datac(\id_inst[13]~q ),
	.datad(\id_inst[4]~q ),
	.cin(gnd),
	.combout(\ex_ctrl_mem_wr~11_combout ),
	.cout());
defparam \ex_ctrl_mem_wr~11 .lut_mask = 16'h001F;
defparam \ex_ctrl_mem_wr~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ex_ctrl_mem_wr~13 (
	.dataa(\id_inst[5]~q ),
	.datab(\id_inst[6]~q ),
	.datac(\ex_ctrl_mem_wr~7_combout ),
	.datad(\ex_ctrl_mem_wr~11_combout ),
	.cin(gnd),
	.combout(\ex_ctrl_mem_wr~13_combout ),
	.cout());
defparam \ex_ctrl_mem_wr~13 .lut_mask = 16'h1000;
defparam \ex_ctrl_mem_wr~13 .sum_lutc_input = "datac";

dffeas \ex_ctrl_mem_wr.01 (
	.clk(clk_clk),
	.d(\ex_ctrl_mem_wr~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\id_pc[7]~31_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\ex_ctrl_mem_wr.01~q ),
	.prn(vcc));
defparam \ex_ctrl_mem_wr.01 .is_wysiwyg = "true";
defparam \ex_ctrl_mem_wr.01 .power_up = "low";

cyclone10lp_lcell_comb \mem_ctrl_mem_wr~10 (
	.dataa(\ex_ctrl_mem_wr.01~q ),
	.datab(\mem_ctrl_mem_wr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_ctrl_mem_wr~10_combout ),
	.cout());
defparam \mem_ctrl_mem_wr~10 .lut_mask = 16'h8888;
defparam \mem_ctrl_mem_wr~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[24]~32 (
	.dataa(data_out_27),
	.datab(mem_rs_1_8),
	.datac(data_out_17),
	.datad(mem_rs_1_16),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[24]~32_combout ),
	.cout());
defparam \io_w_dmem_dat_data[24]~32 .lut_mask = 16'h5E0E;
defparam \io_w_dmem_dat_data[24]~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~66 (
	.dataa(\ex_reg_rs2_bypass[24]~114_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[24]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~66_combout ),
	.cout());
defparam \mem_rs_1~66 .lut_mask = 16'hEA00;
defparam \mem_rs_1~66 .sum_lutc_input = "datac";

dffeas \mem_rs_1[24] (
	.clk(clk_clk),
	.d(\mem_rs_1~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_rs_1[24]~q ),
	.prn(vcc));
defparam \mem_rs_1[24] .is_wysiwyg = "true";
defparam \mem_rs_1[24] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[24]~33 (
	.dataa(mem_rs_1_0),
	.datab(data_out_27),
	.datac(\io_w_dmem_dat_data[24]~32_combout ),
	.datad(\mem_rs_1[24]~q ),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[24]~33_combout ),
	.cout());
defparam \io_w_dmem_dat_data[24]~33 .lut_mask = 16'hF838;
defparam \io_w_dmem_dat_data[24]~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[25]~34 (
	.dataa(data_out_17),
	.datab(mem_rs_1_1),
	.datac(data_out_27),
	.datad(mem_rs_1_17),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[25]~34_combout ),
	.cout());
defparam \io_w_dmem_dat_data[25]~34 .lut_mask = 16'hDAD0;
defparam \io_w_dmem_dat_data[25]~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~67 (
	.dataa(\ex_reg_rs2_bypass[25]~110_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[25]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~67_combout ),
	.cout());
defparam \mem_rs_1~67 .lut_mask = 16'hEA00;
defparam \mem_rs_1~67 .sum_lutc_input = "datac";

dffeas \mem_rs_1[25] (
	.clk(clk_clk),
	.d(\mem_rs_1~67_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_rs_1[25]~q ),
	.prn(vcc));
defparam \mem_rs_1[25] .is_wysiwyg = "true";
defparam \mem_rs_1[25] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[25]~35 (
	.dataa(mem_rs_1_9),
	.datab(data_out_17),
	.datac(\io_w_dmem_dat_data[25]~34_combout ),
	.datad(\mem_rs_1[25]~q ),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[25]~35_combout ),
	.cout());
defparam \io_w_dmem_dat_data[25]~35 .lut_mask = 16'hF2C2;
defparam \io_w_dmem_dat_data[25]~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[26]~36 (
	.dataa(data_out_27),
	.datab(mem_rs_1_10),
	.datac(data_out_17),
	.datad(mem_rs_1_18),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[26]~36_combout ),
	.cout());
defparam \io_w_dmem_dat_data[26]~36 .lut_mask = 16'h5E0E;
defparam \io_w_dmem_dat_data[26]~36 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~68 (
	.dataa(\ex_reg_rs2_bypass[26]~118_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[26]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~68_combout ),
	.cout());
defparam \mem_rs_1~68 .lut_mask = 16'hEA00;
defparam \mem_rs_1~68 .sum_lutc_input = "datac";

dffeas \mem_rs_1[26] (
	.clk(clk_clk),
	.d(\mem_rs_1~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_rs_1[26]~q ),
	.prn(vcc));
defparam \mem_rs_1[26] .is_wysiwyg = "true";
defparam \mem_rs_1[26] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[26]~37 (
	.dataa(mem_rs_1_2),
	.datab(data_out_27),
	.datac(\io_w_dmem_dat_data[26]~36_combout ),
	.datad(\mem_rs_1[26]~q ),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[26]~37_combout ),
	.cout());
defparam \io_w_dmem_dat_data[26]~37 .lut_mask = 16'hF838;
defparam \io_w_dmem_dat_data[26]~37 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[27]~38 (
	.dataa(data_out_17),
	.datab(mem_rs_1_3),
	.datac(data_out_27),
	.datad(mem_rs_1_19),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[27]~38_combout ),
	.cout());
defparam \io_w_dmem_dat_data[27]~38 .lut_mask = 16'hDAD0;
defparam \io_w_dmem_dat_data[27]~38 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~69 (
	.dataa(\ex_reg_rs2_bypass[27]~122_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[27]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~69_combout ),
	.cout());
defparam \mem_rs_1~69 .lut_mask = 16'hEA00;
defparam \mem_rs_1~69 .sum_lutc_input = "datac";

dffeas \mem_rs_1[27] (
	.clk(clk_clk),
	.d(\mem_rs_1~69_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_rs_1[27]~q ),
	.prn(vcc));
defparam \mem_rs_1[27] .is_wysiwyg = "true";
defparam \mem_rs_1[27] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[27]~39 (
	.dataa(mem_rs_1_11),
	.datab(data_out_17),
	.datac(\io_w_dmem_dat_data[27]~38_combout ),
	.datad(\mem_rs_1[27]~q ),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[27]~39_combout ),
	.cout());
defparam \io_w_dmem_dat_data[27]~39 .lut_mask = 16'hF2C2;
defparam \io_w_dmem_dat_data[27]~39 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[28]~40 (
	.dataa(data_out_27),
	.datab(mem_rs_1_12),
	.datac(data_out_17),
	.datad(mem_rs_1_20),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[28]~40_combout ),
	.cout());
defparam \io_w_dmem_dat_data[28]~40 .lut_mask = 16'h5E0E;
defparam \io_w_dmem_dat_data[28]~40 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~70 (
	.dataa(\ex_reg_rs2_bypass[28]~21_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[28]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~70_combout ),
	.cout());
defparam \mem_rs_1~70 .lut_mask = 16'hEA00;
defparam \mem_rs_1~70 .sum_lutc_input = "datac";

dffeas \mem_rs_1[28] (
	.clk(clk_clk),
	.d(\mem_rs_1~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_rs_1[28]~q ),
	.prn(vcc));
defparam \mem_rs_1[28] .is_wysiwyg = "true";
defparam \mem_rs_1[28] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[28]~41 (
	.dataa(mem_rs_1_4),
	.datab(data_out_27),
	.datac(\io_w_dmem_dat_data[28]~40_combout ),
	.datad(\mem_rs_1[28]~q ),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[28]~41_combout ),
	.cout());
defparam \io_w_dmem_dat_data[28]~41 .lut_mask = 16'hF838;
defparam \io_w_dmem_dat_data[28]~41 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[29]~42 (
	.dataa(data_out_17),
	.datab(mem_rs_1_5),
	.datac(data_out_27),
	.datad(mem_rs_1_21),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[29]~42_combout ),
	.cout());
defparam \io_w_dmem_dat_data[29]~42 .lut_mask = 16'hDAD0;
defparam \io_w_dmem_dat_data[29]~42 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~71 (
	.dataa(\ex_reg_rs2_bypass[29]~17_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[29]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~71_combout ),
	.cout());
defparam \mem_rs_1~71 .lut_mask = 16'hEA00;
defparam \mem_rs_1~71 .sum_lutc_input = "datac";

dffeas \mem_rs_1[29] (
	.clk(clk_clk),
	.d(\mem_rs_1~71_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_rs_1[29]~q ),
	.prn(vcc));
defparam \mem_rs_1[29] .is_wysiwyg = "true";
defparam \mem_rs_1[29] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[29]~43 (
	.dataa(mem_rs_1_13),
	.datab(data_out_17),
	.datac(\io_w_dmem_dat_data[29]~42_combout ),
	.datad(\mem_rs_1[29]~q ),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[29]~43_combout ),
	.cout());
defparam \io_w_dmem_dat_data[29]~43 .lut_mask = 16'hF2C2;
defparam \io_w_dmem_dat_data[29]~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[30]~44 (
	.dataa(data_out_27),
	.datab(mem_rs_1_14),
	.datac(data_out_17),
	.datad(mem_rs_1_22),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[30]~44_combout ),
	.cout());
defparam \io_w_dmem_dat_data[30]~44 .lut_mask = 16'h5E0E;
defparam \io_w_dmem_dat_data[30]~44 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~72 (
	.dataa(\ex_reg_rs2_bypass[30]~25_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[30]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~72_combout ),
	.cout());
defparam \mem_rs_1~72 .lut_mask = 16'hEA00;
defparam \mem_rs_1~72 .sum_lutc_input = "datac";

dffeas \mem_rs_1[30] (
	.clk(clk_clk),
	.d(\mem_rs_1~72_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_rs_1[30]~q ),
	.prn(vcc));
defparam \mem_rs_1[30] .is_wysiwyg = "true";
defparam \mem_rs_1[30] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[30]~45 (
	.dataa(mem_rs_1_6),
	.datab(data_out_27),
	.datac(\io_w_dmem_dat_data[30]~44_combout ),
	.datad(\mem_rs_1[30]~q ),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[30]~45_combout ),
	.cout());
defparam \io_w_dmem_dat_data[30]~45 .lut_mask = 16'hF838;
defparam \io_w_dmem_dat_data[30]~45 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[31]~46 (
	.dataa(data_out_17),
	.datab(mem_rs_1_7),
	.datac(data_out_27),
	.datad(mem_rs_1_23),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[31]~46_combout ),
	.cout());
defparam \io_w_dmem_dat_data[31]~46 .lut_mask = 16'hDAD0;
defparam \io_w_dmem_dat_data[31]~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mem_rs_1~73 (
	.dataa(\ex_reg_rs2_bypass[31]~29_combout ),
	.datab(\_T_3681~3_combout ),
	.datac(\mem_csr_data[31]~q ),
	.datad(\mem_ctrl_mem_wr~7_combout ),
	.cin(gnd),
	.combout(\mem_rs_1~73_combout ),
	.cout());
defparam \mem_rs_1~73 .lut_mask = 16'hEA00;
defparam \mem_rs_1~73 .sum_lutc_input = "datac";

dffeas \mem_rs_1[31] (
	.clk(clk_clk),
	.d(\mem_rs_1~73_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_rs_1[31]~q ),
	.prn(vcc));
defparam \mem_rs_1[31] .is_wysiwyg = "true";
defparam \mem_rs_1[31] .power_up = "low";

cyclone10lp_lcell_comb \io_w_dmem_dat_data[31]~47 (
	.dataa(mem_rs_1_15),
	.datab(data_out_17),
	.datac(\io_w_dmem_dat_data[31]~46_combout ),
	.datad(\mem_rs_1[31]~q ),
	.cin(gnd),
	.combout(\io_w_dmem_dat_data[31]~47_combout ),
	.cout());
defparam \io_w_dmem_dat_data[31]~47 .lut_mask = 16'hF2C2;
defparam \io_w_dmem_dat_data[31]~47 .sum_lutc_input = "datac";

endmodule

module kyogenrv_fpga_ALU (
	ex_ctrl_alu_op1_0,
	ex_ctrl_alu_op1_1,
	ex_ctrl_imm_type011,
	ex_ctrl_alu_func_0,
	_T_3_0,
	_T_3_1,
	_T_3_2,
	_T_3_3,
	_T_3_4,
	_T_3_5,
	_T_3_6,
	_T_3_7,
	_T_3_8,
	_T_3_9,
	_T_3_10,
	_T_3_11,
	_T_3_12,
	_T_3_13,
	_T_3_14,
	_T_3_15,
	_T_3_16,
	_T_3_17,
	_T_3_18,
	_T_3_19,
	_T_3_20,
	_T_3_21,
	_T_3_22,
	_T_3_23,
	_T_3_24,
	_T_3_25,
	_T_3_26,
	_T_3_27,
	_T_3_28,
	_T_3_29,
	_T_3_30,
	_T_3_31,
	csr_io_alu_op1_0,
	ex_ctrl_alu_op201,
	ex_ctrl_alu_op210,
	csr_io_alu_op2_1,
	ex_reg_rs2_bypass_1,
	io_sw_r_ex_imm_1,
	csr_io_alu_op2_11,
	csr_io_alu_op2_0,
	alu_io_op2_3,
	ex_reg_rs2_bypass_0,
	_T_3681,
	ex_reg_rs2_bypass_01,
	csr_io_alu_op2_01,
	_T_123_31,
	alu_io_op2_9,
	alu_io_op2_8,
	alu_io_op2_10,
	alu_io_op2_11,
	_T_123_11,
	mem_csr_data_12,
	mem_csr_data_13,
	alu_io_op2_13,
	ex_reg_rs2_bypass_13,
	ex_reg_rs2_bypass_131,
	alu_io_op2_12,
	ex_reg_rs2_bypass_12,
	mem_csr_data_14,
	alu_io_op2_14,
	ex_reg_rs2_bypass_14,
	ex_reg_rs2_bypass_15,
	alu_io_op2_15,
	_T_123_15,
	alu_io_op2_17,
	ex_reg_rs2_bypass_17,
	alu_io_op2_16,
	ex_reg_rs2_bypass_16,
	alu_io_op2_18,
	ex_reg_rs2_bypass_18,
	ex_reg_rs2_bypass_19,
	alu_io_op2_19,
	_T_123_19,
	alu_io_op2_4,
	io_sw_r_ex_imm_4,
	alu_io_op2_41,
	ex_ctrl_alu_func_3,
	alu_io_op2_2,
	_T_123_2,
	alu_io_op2_31,
	io_sw_r_ex_imm_3,
	alu_io_op2_32,
	alu_io_op2_5,
	alu_io_op2_6,
	alu_io_op2_7,
	_T_123_7,
	alu_io_op1_23,
	alu_io_op1_27,
	ex_ctrl_alu_func_1,
	ex_ctrl_alu_func_2,
	LessThan0,
	_T_125,
	alu_io_op1_31,
	csr_io_alu_op1_01,
	alu_io_op1_30,
	csr_io_alu_op1_1,
	ShiftRight0,
	alu_io_op1_8,
	alu_io_op1_7,
	alu_io_op1_24,
	alu_io_op1_4,
	alu_io_op1_3,
	alu_io_op1_28,
	alu_io_op1_6,
	alu_io_op1_25,
	alu_io_op1_5,
	alu_io_op1_26,
	alu_io_op1_2,
	alu_io_op1_29,
	alu_io_op1_12,
	alu_io_op1_19,
	alu_io_op1_11,
	alu_io_op1_20,
	alu_io_op1_10,
	alu_io_op1_21,
	alu_io_op1_9,
	alu_io_op1_22,
	alu_io_op1_16,
	alu_io_op1_15,
	alu_io_op1_14,
	alu_io_op1_17,
	alu_io_op1_13,
	alu_io_op1_18,
	ShiftRight01,
	ShiftRight02,
	ShiftRight03,
	io_out_0,
	ShiftRight04,
	ShiftRight05,
	ShiftRight06,
	ShiftRight07,
	ShiftRight08,
	ShiftRight09,
	ShiftRight010,
	ShiftRight011,
	ShiftRight012,
	ShiftRight013,
	ShiftRight014,
	ShiftRight015,
	ShiftRight016,
	ShiftRight017,
	_T_123_13,
	ShiftRight018,
	ShiftRight019,
	ShiftRight020,
	ShiftRight021,
	_T_139_18,
	ShiftRight022,
	ShiftRight023,
	ShiftRight024,
	ShiftRight025,
	csr_io_alu_op1_11,
	csr_io_alu_op1_02,
	alu_io_op1_281,
	alu_io_op1_291,
	alu_io_op2_29,
	alu_io_op2_28,
	alu_io_op1_301,
	alu_io_op2_30,
	alu_io_op1_311,
	alu_io_op2_311,
	alu_io_op1_81,
	alu_io_op1_91,
	alu_io_op1_101,
	alu_io_op1_111,
	alu_io_op1_121,
	alu_io_op1_131,
	alu_io_op2_131,
	alu_io_op2_121,
	alu_io_op1_141,
	alu_io_op2_141,
	alu_io_op1_151,
	alu_io_op1_161,
	alu_io_op1_171,
	alu_io_op2_171,
	alu_io_op2_161,
	alu_io_op1_181,
	alu_io_op2_181,
	alu_io_op1_191,
	alu_io_op1_41,
	alu_io_op1_210,
	alu_io_op1_51,
	alu_io_op1_32,
	alu_io_op1_61,
	alu_io_op1_71,
	alu_io_op1_201,
	alu_io_op1_211,
	alu_io_op2_21,
	alu_io_op2_20,
	alu_io_op1_221,
	alu_io_op2_22,
	alu_io_op2_23,
	_T_123_23,
	alu_io_op1_241,
	alu_io_op1_251,
	alu_io_op2_25,
	alu_io_op2_24,
	alu_io_op1_261,
	alu_io_op2_26,
	alu_io_op2_27,
	_T_123_27,
	alu_io_op1_271,
	alu_io_op1_231,
	alu_io_op2_210,
	_T_123_29,
	ShiftRight026,
	ShiftRight027,
	_T_123_17,
	ShiftRight028,
	ShiftRight029,
	ShiftRight030,
	ShiftRight031,
	_T_123_21,
	_T_123_25)/* synthesis synthesis_greybox=0 */;
input 	ex_ctrl_alu_op1_0;
input 	ex_ctrl_alu_op1_1;
input 	ex_ctrl_imm_type011;
input 	ex_ctrl_alu_func_0;
output 	_T_3_0;
output 	_T_3_1;
output 	_T_3_2;
output 	_T_3_3;
output 	_T_3_4;
output 	_T_3_5;
output 	_T_3_6;
output 	_T_3_7;
output 	_T_3_8;
output 	_T_3_9;
output 	_T_3_10;
output 	_T_3_11;
output 	_T_3_12;
output 	_T_3_13;
output 	_T_3_14;
output 	_T_3_15;
output 	_T_3_16;
output 	_T_3_17;
output 	_T_3_18;
output 	_T_3_19;
output 	_T_3_20;
output 	_T_3_21;
output 	_T_3_22;
output 	_T_3_23;
output 	_T_3_24;
output 	_T_3_25;
output 	_T_3_26;
output 	_T_3_27;
output 	_T_3_28;
output 	_T_3_29;
output 	_T_3_30;
output 	_T_3_31;
input 	csr_io_alu_op1_0;
input 	ex_ctrl_alu_op201;
input 	ex_ctrl_alu_op210;
input 	csr_io_alu_op2_1;
input 	ex_reg_rs2_bypass_1;
input 	io_sw_r_ex_imm_1;
input 	csr_io_alu_op2_11;
input 	csr_io_alu_op2_0;
input 	alu_io_op2_3;
input 	ex_reg_rs2_bypass_0;
input 	_T_3681;
input 	ex_reg_rs2_bypass_01;
input 	csr_io_alu_op2_01;
output 	_T_123_31;
input 	alu_io_op2_9;
input 	alu_io_op2_8;
input 	alu_io_op2_10;
input 	alu_io_op2_11;
output 	_T_123_11;
input 	mem_csr_data_12;
input 	mem_csr_data_13;
input 	alu_io_op2_13;
input 	ex_reg_rs2_bypass_13;
input 	ex_reg_rs2_bypass_131;
input 	alu_io_op2_12;
input 	ex_reg_rs2_bypass_12;
input 	mem_csr_data_14;
input 	alu_io_op2_14;
input 	ex_reg_rs2_bypass_14;
input 	ex_reg_rs2_bypass_15;
input 	alu_io_op2_15;
output 	_T_123_15;
input 	alu_io_op2_17;
input 	ex_reg_rs2_bypass_17;
input 	alu_io_op2_16;
input 	ex_reg_rs2_bypass_16;
input 	alu_io_op2_18;
input 	ex_reg_rs2_bypass_18;
input 	ex_reg_rs2_bypass_19;
input 	alu_io_op2_19;
output 	_T_123_19;
input 	alu_io_op2_4;
input 	io_sw_r_ex_imm_4;
input 	alu_io_op2_41;
input 	ex_ctrl_alu_func_3;
input 	alu_io_op2_2;
output 	_T_123_2;
input 	alu_io_op2_31;
input 	io_sw_r_ex_imm_3;
input 	alu_io_op2_32;
input 	alu_io_op2_5;
input 	alu_io_op2_6;
input 	alu_io_op2_7;
output 	_T_123_7;
input 	alu_io_op1_23;
input 	alu_io_op1_27;
input 	ex_ctrl_alu_func_1;
input 	ex_ctrl_alu_func_2;
output 	LessThan0;
output 	_T_125;
input 	alu_io_op1_31;
input 	csr_io_alu_op1_01;
input 	alu_io_op1_30;
input 	csr_io_alu_op1_1;
output 	ShiftRight0;
input 	alu_io_op1_8;
input 	alu_io_op1_7;
input 	alu_io_op1_24;
input 	alu_io_op1_4;
input 	alu_io_op1_3;
input 	alu_io_op1_28;
input 	alu_io_op1_6;
input 	alu_io_op1_25;
input 	alu_io_op1_5;
input 	alu_io_op1_26;
input 	alu_io_op1_2;
input 	alu_io_op1_29;
input 	alu_io_op1_12;
input 	alu_io_op1_19;
input 	alu_io_op1_11;
input 	alu_io_op1_20;
input 	alu_io_op1_10;
input 	alu_io_op1_21;
input 	alu_io_op1_9;
input 	alu_io_op1_22;
input 	alu_io_op1_16;
input 	alu_io_op1_15;
input 	alu_io_op1_14;
input 	alu_io_op1_17;
input 	alu_io_op1_13;
input 	alu_io_op1_18;
output 	ShiftRight01;
output 	ShiftRight02;
output 	ShiftRight03;
output 	io_out_0;
output 	ShiftRight04;
output 	ShiftRight05;
output 	ShiftRight06;
output 	ShiftRight07;
output 	ShiftRight08;
output 	ShiftRight09;
output 	ShiftRight010;
output 	ShiftRight011;
output 	ShiftRight012;
output 	ShiftRight013;
output 	ShiftRight014;
output 	ShiftRight015;
output 	ShiftRight016;
output 	ShiftRight017;
output 	_T_123_13;
output 	ShiftRight018;
output 	ShiftRight019;
output 	ShiftRight020;
output 	ShiftRight021;
output 	_T_139_18;
output 	ShiftRight022;
output 	ShiftRight023;
output 	ShiftRight024;
output 	ShiftRight025;
input 	csr_io_alu_op1_11;
input 	csr_io_alu_op1_02;
input 	alu_io_op1_281;
input 	alu_io_op1_291;
input 	alu_io_op2_29;
input 	alu_io_op2_28;
input 	alu_io_op1_301;
input 	alu_io_op2_30;
input 	alu_io_op1_311;
input 	alu_io_op2_311;
input 	alu_io_op1_81;
input 	alu_io_op1_91;
input 	alu_io_op1_101;
input 	alu_io_op1_111;
input 	alu_io_op1_121;
input 	alu_io_op1_131;
input 	alu_io_op2_131;
input 	alu_io_op2_121;
input 	alu_io_op1_141;
input 	alu_io_op2_141;
input 	alu_io_op1_151;
input 	alu_io_op1_161;
input 	alu_io_op1_171;
input 	alu_io_op2_171;
input 	alu_io_op2_161;
input 	alu_io_op1_181;
input 	alu_io_op2_181;
input 	alu_io_op1_191;
input 	alu_io_op1_41;
input 	alu_io_op1_210;
input 	alu_io_op1_51;
input 	alu_io_op1_32;
input 	alu_io_op1_61;
input 	alu_io_op1_71;
input 	alu_io_op1_201;
input 	alu_io_op1_211;
input 	alu_io_op2_21;
input 	alu_io_op2_20;
input 	alu_io_op1_221;
input 	alu_io_op2_22;
input 	alu_io_op2_23;
output 	_T_123_23;
input 	alu_io_op1_241;
input 	alu_io_op1_251;
input 	alu_io_op2_25;
input 	alu_io_op2_24;
input 	alu_io_op1_261;
input 	alu_io_op2_26;
input 	alu_io_op2_27;
output 	_T_123_27;
input 	alu_io_op1_271;
input 	alu_io_op1_231;
input 	alu_io_op2_210;
output 	_T_123_29;
output 	ShiftRight026;
output 	ShiftRight027;
output 	_T_123_17;
output 	ShiftRight028;
output 	ShiftRight029;
output 	ShiftRight030;
output 	ShiftRight031;
output 	_T_123_21;
output 	_T_123_25;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_T_3[0]~1 ;
wire \_T_3[1]~3 ;
wire \_T_3[2]~5 ;
wire \_T_3[3]~7 ;
wire \_T_3[4]~9 ;
wire \_T_3[5]~11 ;
wire \_T_3[6]~13 ;
wire \_T_3[7]~15 ;
wire \_T_3[8]~17 ;
wire \_T_3[9]~19 ;
wire \_T_3[10]~21 ;
wire \_T_3[11]~23 ;
wire \_T_3[12]~25 ;
wire \_T_3[13]~27 ;
wire \_T_3[14]~29 ;
wire \_T_3[15]~31 ;
wire \_T_3[16]~33 ;
wire \_T_3[17]~35 ;
wire \_T_3[18]~37 ;
wire \_T_3[19]~39 ;
wire \_T_3[20]~41 ;
wire \_T_3[21]~43 ;
wire \_T_3[22]~45 ;
wire \_T_3[23]~47 ;
wire \_T_3[24]~49 ;
wire \_T_3[25]~51 ;
wire \_T_3[26]~53 ;
wire \_T_3[27]~55 ;
wire \_T_3[28]~57 ;
wire \_T_3[29]~59 ;
wire \_T_3[30]~61 ;
wire \op2_inv[0]~46_combout ;
wire \op2_inv[0]~42_combout ;
wire \Add0~1_cout ;
wire \op2_inv[1]~45_combout ;
wire \op2_inv[1]~41_combout ;
wire \op2_inv[2]~40_combout ;
wire \op2_inv[3]~38_combout ;
wire \op2_inv[3]~39_combout ;
wire \op2_inv[4]~36_combout ;
wire \op2_inv[4]~37_combout ;
wire \op2_inv[5]~35_combout ;
wire \op2_inv[6]~34_combout ;
wire \op2_inv[7]~33_combout ;
wire \op2_inv[8]~32_combout ;
wire \op2_inv[9]~31_combout ;
wire \op2_inv[10]~30_combout ;
wire \op2_inv[11]~29_combout ;
wire \op2_inv[12]~27_combout ;
wire \op2_inv[12]~28_combout ;
wire \op2_inv[13]~25_combout ;
wire \op2_inv[13]~26_combout ;
wire \op2_inv[14]~23_combout ;
wire \op2_inv[14]~24_combout ;
wire \op2_inv[15]~22_combout ;
wire \op2_inv[16]~21_combout ;
wire \op2_inv[17]~20_combout ;
wire \op2_inv[18]~19_combout ;
wire \op2_inv[19]~18_combout ;
wire \op2_inv[20]~17_combout ;
wire \op2_inv[21]~16_combout ;
wire \op2_inv[22]~15_combout ;
wire \op2_inv[23]~14_combout ;
wire \op2_inv[24]~13_combout ;
wire \op2_inv[25]~12_combout ;
wire \op2_inv[26]~11_combout ;
wire \op2_inv[27]~10_combout ;
wire \op2_inv[28]~9_combout ;
wire \op2_inv[29]~8_combout ;
wire \op2_inv[30]~7_combout ;
wire \op2_inv[31]~6_combout ;
wire \_T_125~0_combout ;
wire \_T_125~1_combout ;
wire \_T_125~2_combout ;
wire \_T_125~3_combout ;
wire \_T_125~4_combout ;
wire \_T_125~5_combout ;
wire \_T_125~6_combout ;
wire \_T_125~7_combout ;
wire \_T_125~8_combout ;
wire \_T_125~9_combout ;
wire \_T_125~10_combout ;
wire \_T_125~11_combout ;
wire \_T_125~12_combout ;
wire \_T_125~13_combout ;
wire \_T_125~14_combout ;
wire \_T_125~15_combout ;
wire \_T_125~16_combout ;
wire \_T_125~17_combout ;
wire \_T_125~18_combout ;
wire \_T_125~19_combout ;
wire \ShiftRight0~241_combout ;
wire \_T_8~0_combout ;
wire \ShiftRight0~32_combout ;
wire \ShiftRight0~33_combout ;
wire \ShiftRight0~34_combout ;
wire \ShiftRight0~35_combout ;
wire \ShiftRight0~242_combout ;
wire \ShiftRight0~36_combout ;
wire \_T_60~combout ;
wire \ShiftRight0~37_combout ;
wire \ShiftRight0~39_combout ;
wire \ShiftRight0~40_combout ;
wire \ShiftRight0~41_combout ;
wire \ShiftRight0~42_combout ;
wire \ShiftRight0~43_combout ;
wire \ShiftRight0~44_combout ;
wire \ShiftRight0~45_combout ;
wire \ShiftRight0~46_combout ;
wire \ShiftRight0~47_combout ;
wire \ShiftRight0~48_combout ;
wire \ShiftRight0~49_combout ;
wire \ShiftRight0~50_combout ;
wire \ShiftRight0~51_combout ;
wire \ShiftRight0~52_combout ;
wire \ShiftRight0~53_combout ;
wire \ShiftRight0~54_combout ;
wire \ShiftRight0~55_combout ;
wire \ShiftRight0~56_combout ;
wire \ShiftRight0~57_combout ;
wire \ShiftRight0~58_combout ;
wire \ShiftRight0~59_combout ;
wire \ShiftRight0~60_combout ;
wire \ShiftRight0~61_combout ;
wire \ShiftRight0~62_combout ;
wire \ShiftRight0~63_combout ;
wire \ShiftRight0~64_combout ;
wire \ShiftRight0~65_combout ;
wire \ShiftRight0~66_combout ;
wire \_T_62[31]~0_combout ;
wire \ShiftRight0~67_combout ;
wire \ShiftRight0~68_combout ;
wire \ShiftRight0~69_combout ;
wire \ShiftRight0~70_combout ;
wire \ShiftRight0~71_combout ;
wire \ShiftRight0~72_combout ;
wire \ShiftRight0~73_combout ;
wire \ShiftRight0~74_combout ;
wire \ShiftRight0~75_combout ;
wire \ShiftRight0~76_combout ;
wire \ShiftRight0~77_combout ;
wire \ShiftRight0~78_combout ;
wire \ShiftRight0~79_combout ;
wire \ShiftRight0~80_combout ;
wire \ShiftRight0~81_combout ;
wire \ShiftRight0~82_combout ;
wire \ShiftRight0~83_combout ;
wire \ShiftRight0~84_combout ;
wire \ShiftRight0~85_combout ;
wire \ShiftRight0~86_combout ;
wire \ShiftRight0~87_combout ;
wire \ShiftRight0~88_combout ;
wire \ShiftRight0~89_combout ;
wire \ShiftRight0~90_combout ;
wire \ShiftRight0~91_combout ;
wire \ShiftRight0~92_combout ;
wire \ShiftRight0~243_combout ;
wire \ShiftRight0~93_combout ;
wire \ShiftRight0~95_combout ;
wire \ShiftRight0~96_combout ;
wire \ShiftRight0~97_combout ;
wire \ShiftRight0~98_combout ;
wire \ShiftRight0~99_combout ;
wire \ShiftRight0~100_combout ;
wire \ShiftRight0~101_combout ;
wire \ShiftRight0~102_combout ;
wire \ShiftRight0~103_combout ;
wire \ShiftRight0~104_combout ;
wire \ShiftRight0~105_combout ;
wire \ShiftRight0~106_combout ;
wire \ShiftRight0~107_combout ;
wire \ShiftRight0~108_combout ;
wire \ShiftRight0~109_combout ;
wire \ShiftRight0~110_combout ;
wire \ShiftRight0~111_combout ;
wire \ShiftRight0~112_combout ;
wire \ShiftRight0~113_combout ;
wire \ShiftRight0~114_combout ;
wire \ShiftRight0~115_combout ;
wire \ShiftRight0~116_combout ;
wire \ShiftRight0~117_combout ;
wire \ShiftRight0~118_combout ;
wire \ShiftRight0~119_combout ;
wire \ShiftRight0~120_combout ;
wire \ShiftRight0~121_combout ;
wire \ShiftRight0~122_combout ;
wire \ShiftRight0~123_combout ;
wire \ShiftRight0~124_combout ;
wire \ShiftRight0~125_combout ;
wire \ShiftRight0~127_combout ;
wire \op2_inv[31]~47_combout ;
wire \op2_inv[31]~43_combout ;
wire \io_out[0]~0_combout ;
wire \op2_inv[31]~44_combout ;
wire \ShiftRight0~129_combout ;
wire \ShiftRight0~131_combout ;
wire \ShiftRight0~132_combout ;
wire \ShiftRight0~133_combout ;
wire \ShiftRight0~134_combout ;
wire \ShiftRight0~135_combout ;
wire \ShiftRight0~136_combout ;
wire \ShiftRight0~137_combout ;
wire \ShiftRight0~138_combout ;
wire \ShiftRight0~139_combout ;
wire \ShiftRight0~140_combout ;
wire \ShiftRight0~141_combout ;
wire \ShiftRight0~142_combout ;
wire \ShiftRight0~143_combout ;
wire \ShiftRight0~144_combout ;
wire \ShiftRight0~145_combout ;
wire \ShiftRight0~146_combout ;
wire \ShiftRight0~147_combout ;
wire \ShiftRight0~148_combout ;
wire \ShiftRight0~149_combout ;
wire \ShiftRight0~151_combout ;
wire \ShiftRight0~153_combout ;
wire \ShiftRight0~154_combout ;
wire \ShiftRight0~155_combout ;
wire \ShiftRight0~156_combout ;
wire \ShiftRight0~157_combout ;
wire \ShiftRight0~244_combout ;
wire \ShiftRight0~158_combout ;
wire \ShiftRight0~159_combout ;
wire \ShiftRight0~160_combout ;
wire \ShiftRight0~161_combout ;
wire \ShiftRight0~162_combout ;
wire \ShiftRight0~163_combout ;
wire \ShiftRight0~164_combout ;
wire \ShiftRight0~165_combout ;
wire \ShiftRight0~166_combout ;
wire \ShiftRight0~168_combout ;
wire \ShiftRight0~169_combout ;
wire \ShiftRight0~170_combout ;
wire \ShiftRight0~171_combout ;
wire \ShiftRight0~172_combout ;
wire \ShiftRight0~245_combout ;
wire \ShiftRight0~246_combout ;
wire \ShiftRight0~247_combout ;
wire \ShiftRight0~174_combout ;
wire \ShiftRight0~176_combout ;
wire \ShiftRight0~177_combout ;
wire \ShiftRight0~178_combout ;
wire \ShiftRight0~179_combout ;
wire \ShiftRight0~181_combout ;
wire \ShiftRight0~182_combout ;
wire \ShiftRight0~184_combout ;
wire \ShiftRight0~185_combout ;
wire \ShiftRight0~186_combout ;
wire \ShiftRight0~187_combout ;
wire \ShiftRight0~189_combout ;
wire \ShiftRight0~191_combout ;
wire \ShiftRight0~192_combout ;
wire \ShiftRight0~193_combout ;
wire \ShiftRight0~194_combout ;
wire \ShiftRight0~196_combout ;
wire \ShiftRight0~248_combout ;
wire \ShiftRight0~199_combout ;
wire \ShiftRight0~200_combout ;
wire \ShiftRight0~201_combout ;
wire \ShiftRight0~202_combout ;
wire \ShiftRight0~205_combout ;
wire \ShiftRight0~206_combout ;
wire \ShiftRight0~207_combout ;
wire \ShiftRight0~208_combout ;
wire \ShiftRight0~211_combout ;
wire \ShiftRight0~212_combout ;
wire \ShiftRight0~213_combout ;
wire \ShiftRight0~214_combout ;
wire \ShiftRight0~215_combout ;
wire \ShiftRight0~218_combout ;
wire \ShiftRight0~219_combout ;
wire \ShiftRight0~220_combout ;
wire \ShiftRight0~221_combout ;
wire \ShiftRight0~223_combout ;
wire \ShiftRight0~224_combout ;
wire \ShiftRight0~225_combout ;
wire \ShiftRight0~252_combout ;
wire \ShiftRight0~226_combout ;
wire \ShiftRight0~227_combout ;
wire \ShiftRight0~229_combout ;
wire \ShiftRight0~230_combout ;
wire \ShiftRight0~231_combout ;
wire \ShiftRight0~232_combout ;
wire \ShiftRight0~234_combout ;
wire \ShiftRight0~255_combout ;
wire \ShiftRight0~235_combout ;
wire \ShiftRight0~237_combout ;
wire \ShiftRight0~238_combout ;
wire \ShiftRight0~239_combout ;
wire \ShiftRight0~204_combout ;
wire \ShiftRight0~210_combout ;


cyclone10lp_lcell_comb \_T_3[0]~0 (
	.dataa(csr_io_alu_op1_02),
	.datab(\op2_inv[0]~42_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1_cout ),
	.combout(_T_3_0),
	.cout(\_T_3[0]~1 ));
defparam \_T_3[0]~0 .lut_mask = 16'h9617;
defparam \_T_3[0]~0 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[1]~2 (
	.dataa(csr_io_alu_op1_11),
	.datab(\op2_inv[1]~41_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[0]~1 ),
	.combout(_T_3_1),
	.cout(\_T_3[1]~3 ));
defparam \_T_3[1]~2 .lut_mask = 16'h698E;
defparam \_T_3[1]~2 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[2]~4 (
	.dataa(alu_io_op1_210),
	.datab(\op2_inv[2]~40_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[1]~3 ),
	.combout(_T_3_2),
	.cout(\_T_3[2]~5 ));
defparam \_T_3[2]~4 .lut_mask = 16'h9617;
defparam \_T_3[2]~4 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[3]~6 (
	.dataa(alu_io_op1_32),
	.datab(\op2_inv[3]~39_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[2]~5 ),
	.combout(_T_3_3),
	.cout(\_T_3[3]~7 ));
defparam \_T_3[3]~6 .lut_mask = 16'h698E;
defparam \_T_3[3]~6 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[4]~8 (
	.dataa(alu_io_op1_41),
	.datab(\op2_inv[4]~37_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[3]~7 ),
	.combout(_T_3_4),
	.cout(\_T_3[4]~9 ));
defparam \_T_3[4]~8 .lut_mask = 16'h9617;
defparam \_T_3[4]~8 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[5]~10 (
	.dataa(alu_io_op1_51),
	.datab(\op2_inv[5]~35_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[4]~9 ),
	.combout(_T_3_5),
	.cout(\_T_3[5]~11 ));
defparam \_T_3[5]~10 .lut_mask = 16'h698E;
defparam \_T_3[5]~10 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[6]~12 (
	.dataa(alu_io_op1_61),
	.datab(\op2_inv[6]~34_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[5]~11 ),
	.combout(_T_3_6),
	.cout(\_T_3[6]~13 ));
defparam \_T_3[6]~12 .lut_mask = 16'h9617;
defparam \_T_3[6]~12 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[7]~14 (
	.dataa(alu_io_op1_71),
	.datab(\op2_inv[7]~33_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[6]~13 ),
	.combout(_T_3_7),
	.cout(\_T_3[7]~15 ));
defparam \_T_3[7]~14 .lut_mask = 16'h698E;
defparam \_T_3[7]~14 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[8]~16 (
	.dataa(alu_io_op1_81),
	.datab(\op2_inv[8]~32_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[7]~15 ),
	.combout(_T_3_8),
	.cout(\_T_3[8]~17 ));
defparam \_T_3[8]~16 .lut_mask = 16'h9617;
defparam \_T_3[8]~16 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[9]~18 (
	.dataa(alu_io_op1_91),
	.datab(\op2_inv[9]~31_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[8]~17 ),
	.combout(_T_3_9),
	.cout(\_T_3[9]~19 ));
defparam \_T_3[9]~18 .lut_mask = 16'h698E;
defparam \_T_3[9]~18 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[10]~20 (
	.dataa(alu_io_op1_101),
	.datab(\op2_inv[10]~30_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[9]~19 ),
	.combout(_T_3_10),
	.cout(\_T_3[10]~21 ));
defparam \_T_3[10]~20 .lut_mask = 16'h9617;
defparam \_T_3[10]~20 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[11]~22 (
	.dataa(alu_io_op1_111),
	.datab(\op2_inv[11]~29_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[10]~21 ),
	.combout(_T_3_11),
	.cout(\_T_3[11]~23 ));
defparam \_T_3[11]~22 .lut_mask = 16'h698E;
defparam \_T_3[11]~22 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[12]~24 (
	.dataa(alu_io_op1_121),
	.datab(\op2_inv[12]~28_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[11]~23 ),
	.combout(_T_3_12),
	.cout(\_T_3[12]~25 ));
defparam \_T_3[12]~24 .lut_mask = 16'h9617;
defparam \_T_3[12]~24 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[13]~26 (
	.dataa(alu_io_op1_131),
	.datab(\op2_inv[13]~26_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[12]~25 ),
	.combout(_T_3_13),
	.cout(\_T_3[13]~27 ));
defparam \_T_3[13]~26 .lut_mask = 16'h698E;
defparam \_T_3[13]~26 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[14]~28 (
	.dataa(alu_io_op1_141),
	.datab(\op2_inv[14]~24_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[13]~27 ),
	.combout(_T_3_14),
	.cout(\_T_3[14]~29 ));
defparam \_T_3[14]~28 .lut_mask = 16'h9617;
defparam \_T_3[14]~28 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[15]~30 (
	.dataa(alu_io_op1_151),
	.datab(\op2_inv[15]~22_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[14]~29 ),
	.combout(_T_3_15),
	.cout(\_T_3[15]~31 ));
defparam \_T_3[15]~30 .lut_mask = 16'h698E;
defparam \_T_3[15]~30 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[16]~32 (
	.dataa(alu_io_op1_161),
	.datab(\op2_inv[16]~21_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[15]~31 ),
	.combout(_T_3_16),
	.cout(\_T_3[16]~33 ));
defparam \_T_3[16]~32 .lut_mask = 16'h9617;
defparam \_T_3[16]~32 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[17]~34 (
	.dataa(alu_io_op1_171),
	.datab(\op2_inv[17]~20_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[16]~33 ),
	.combout(_T_3_17),
	.cout(\_T_3[17]~35 ));
defparam \_T_3[17]~34 .lut_mask = 16'h698E;
defparam \_T_3[17]~34 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[18]~36 (
	.dataa(alu_io_op1_181),
	.datab(\op2_inv[18]~19_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[17]~35 ),
	.combout(_T_3_18),
	.cout(\_T_3[18]~37 ));
defparam \_T_3[18]~36 .lut_mask = 16'h9617;
defparam \_T_3[18]~36 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[19]~38 (
	.dataa(alu_io_op1_191),
	.datab(\op2_inv[19]~18_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[18]~37 ),
	.combout(_T_3_19),
	.cout(\_T_3[19]~39 ));
defparam \_T_3[19]~38 .lut_mask = 16'h698E;
defparam \_T_3[19]~38 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[20]~40 (
	.dataa(alu_io_op1_201),
	.datab(\op2_inv[20]~17_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[19]~39 ),
	.combout(_T_3_20),
	.cout(\_T_3[20]~41 ));
defparam \_T_3[20]~40 .lut_mask = 16'h9617;
defparam \_T_3[20]~40 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[21]~42 (
	.dataa(alu_io_op1_211),
	.datab(\op2_inv[21]~16_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[20]~41 ),
	.combout(_T_3_21),
	.cout(\_T_3[21]~43 ));
defparam \_T_3[21]~42 .lut_mask = 16'h698E;
defparam \_T_3[21]~42 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[22]~44 (
	.dataa(alu_io_op1_221),
	.datab(\op2_inv[22]~15_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[21]~43 ),
	.combout(_T_3_22),
	.cout(\_T_3[22]~45 ));
defparam \_T_3[22]~44 .lut_mask = 16'h9617;
defparam \_T_3[22]~44 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[23]~46 (
	.dataa(alu_io_op1_231),
	.datab(\op2_inv[23]~14_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[22]~45 ),
	.combout(_T_3_23),
	.cout(\_T_3[23]~47 ));
defparam \_T_3[23]~46 .lut_mask = 16'h698E;
defparam \_T_3[23]~46 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[24]~48 (
	.dataa(alu_io_op1_241),
	.datab(\op2_inv[24]~13_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[23]~47 ),
	.combout(_T_3_24),
	.cout(\_T_3[24]~49 ));
defparam \_T_3[24]~48 .lut_mask = 16'h9617;
defparam \_T_3[24]~48 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[25]~50 (
	.dataa(alu_io_op1_251),
	.datab(\op2_inv[25]~12_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[24]~49 ),
	.combout(_T_3_25),
	.cout(\_T_3[25]~51 ));
defparam \_T_3[25]~50 .lut_mask = 16'h698E;
defparam \_T_3[25]~50 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[26]~52 (
	.dataa(alu_io_op1_261),
	.datab(\op2_inv[26]~11_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[25]~51 ),
	.combout(_T_3_26),
	.cout(\_T_3[26]~53 ));
defparam \_T_3[26]~52 .lut_mask = 16'h9617;
defparam \_T_3[26]~52 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[27]~54 (
	.dataa(alu_io_op1_271),
	.datab(\op2_inv[27]~10_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[26]~53 ),
	.combout(_T_3_27),
	.cout(\_T_3[27]~55 ));
defparam \_T_3[27]~54 .lut_mask = 16'h698E;
defparam \_T_3[27]~54 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[28]~56 (
	.dataa(alu_io_op1_281),
	.datab(\op2_inv[28]~9_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[27]~55 ),
	.combout(_T_3_28),
	.cout(\_T_3[28]~57 ));
defparam \_T_3[28]~56 .lut_mask = 16'h9617;
defparam \_T_3[28]~56 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[29]~58 (
	.dataa(alu_io_op1_291),
	.datab(\op2_inv[29]~8_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[28]~57 ),
	.combout(_T_3_29),
	.cout(\_T_3[29]~59 ));
defparam \_T_3[29]~58 .lut_mask = 16'h698E;
defparam \_T_3[29]~58 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[30]~60 (
	.dataa(alu_io_op1_301),
	.datab(\op2_inv[30]~7_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\_T_3[29]~59 ),
	.combout(_T_3_30),
	.cout(\_T_3[30]~61 ));
defparam \_T_3[30]~60 .lut_mask = 16'h9617;
defparam \_T_3[30]~60 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_3[31]~62 (
	.dataa(alu_io_op1_311),
	.datab(\op2_inv[31]~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(\_T_3[30]~61 ),
	.combout(_T_3_31),
	.cout());
defparam \_T_3[31]~62 .lut_mask = 16'h6969;
defparam \_T_3[31]~62 .sum_lutc_input = "cin";

cyclone10lp_lcell_comb \_T_123[31] (
	.dataa(gnd),
	.datab(gnd),
	.datac(alu_io_op1_311),
	.datad(alu_io_op2_311),
	.cin(gnd),
	.combout(_T_123_31),
	.cout());
defparam \_T_123[31] .lut_mask = 16'h0FF0;
defparam \_T_123[31] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_123[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(alu_io_op1_111),
	.datad(alu_io_op2_11),
	.cin(gnd),
	.combout(_T_123_11),
	.cout());
defparam \_T_123[11] .lut_mask = 16'h0FF0;
defparam \_T_123[11] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_123[15] (
	.dataa(alu_io_op2_3),
	.datab(ex_reg_rs2_bypass_15),
	.datac(alu_io_op2_15),
	.datad(alu_io_op1_151),
	.cin(gnd),
	.combout(_T_123_15),
	.cout());
defparam \_T_123[15] .lut_mask = 16'h07F8;
defparam \_T_123[15] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_123[19] (
	.dataa(alu_io_op2_3),
	.datab(ex_reg_rs2_bypass_19),
	.datac(alu_io_op2_19),
	.datad(alu_io_op1_191),
	.cin(gnd),
	.combout(_T_123_19),
	.cout());
defparam \_T_123[19] .lut_mask = 16'h07F8;
defparam \_T_123[19] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_123[2] (
	.dataa(gnd),
	.datab(alu_io_op1_210),
	.datac(csr_io_alu_op2_1),
	.datad(alu_io_op2_2),
	.cin(gnd),
	.combout(_T_123_2),
	.cout());
defparam \_T_123[2] .lut_mask = 16'h3CCC;
defparam \_T_123[2] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_123[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(alu_io_op1_71),
	.datad(alu_io_op2_7),
	.cin(gnd),
	.combout(_T_123_7),
	.cout());
defparam \_T_123[7] .lut_mask = 16'h0FF0;
defparam \_T_123[7] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \LessThan0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_1),
	.datad(ex_ctrl_alu_func_2),
	.cin(gnd),
	.combout(LessThan0),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'h0FFF;
defparam \LessThan0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~20 (
	.dataa(\_T_125~1_combout ),
	.datab(\_T_125~9_combout ),
	.datac(\_T_125~17_combout ),
	.datad(\_T_125~19_combout ),
	.cin(gnd),
	.combout(_T_125),
	.cout());
defparam \_T_125~20 .lut_mask = 16'hFF80;
defparam \_T_125~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~38 (
	.dataa(\ShiftRight0~36_combout ),
	.datab(\_T_60~combout ),
	.datac(\ShiftRight0~242_combout ),
	.datad(\ShiftRight0~37_combout ),
	.cin(gnd),
	.combout(ShiftRight0),
	.cout());
defparam \ShiftRight0~38 .lut_mask = 16'hEAEE;
defparam \ShiftRight0~38 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~94 (
	.dataa(\ShiftRight0~66_combout ),
	.datab(\ShiftRight0~93_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(ShiftRight01),
	.cout());
defparam \ShiftRight0~94 .lut_mask = 16'hEEEE;
defparam \ShiftRight0~94 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~126 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~108_combout ),
	.datac(\ShiftRight0~125_combout ),
	.datad(alu_io_op2_41),
	.cin(gnd),
	.combout(ShiftRight02),
	.cout());
defparam \ShiftRight0~126 .lut_mask = 16'h88A0;
defparam \ShiftRight0~126 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~128 (
	.dataa(\_T_60~combout ),
	.datab(\_T_62[31]~0_combout ),
	.datac(alu_io_op2_41),
	.datad(\ShiftRight0~127_combout ),
	.cin(gnd),
	.combout(ShiftRight03),
	.cout());
defparam \ShiftRight0~128 .lut_mask = 16'hAAAC;
defparam \ShiftRight0~128 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[0]~1 (
	.dataa(csr_io_alu_op2_01),
	.datab(ex_ctrl_alu_func_1),
	.datac(\io_out[0]~0_combout ),
	.datad(\op2_inv[31]~44_combout ),
	.cin(gnd),
	.combout(io_out_0),
	.cout());
defparam \io_out[0]~1 .lut_mask = 16'hF838;
defparam \io_out[0]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~130 (
	.dataa(\_T_60~combout ),
	.datab(\ShiftRight0~70_combout ),
	.datac(alu_io_op2_41),
	.datad(\ShiftRight0~129_combout ),
	.cin(gnd),
	.combout(ShiftRight04),
	.cout());
defparam \ShiftRight0~130 .lut_mask = 16'hAAAC;
defparam \ShiftRight0~130 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~150 (
	.dataa(\ShiftRight0~140_combout ),
	.datab(\ShiftRight0~149_combout ),
	.datac(gnd),
	.datad(alu_io_op2_41),
	.cin(gnd),
	.combout(ShiftRight05),
	.cout());
defparam \ShiftRight0~150 .lut_mask = 16'hAAEE;
defparam \ShiftRight0~150 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~152 (
	.dataa(\_T_60~combout ),
	.datab(\ShiftRight0~151_combout ),
	.datac(alu_io_op2_41),
	.datad(\ShiftRight0~129_combout ),
	.cin(gnd),
	.combout(ShiftRight06),
	.cout());
defparam \ShiftRight0~152 .lut_mask = 16'hAAAC;
defparam \ShiftRight0~152 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~167 (
	.dataa(\ShiftRight0~158_combout ),
	.datab(\ShiftRight0~166_combout ),
	.datac(gnd),
	.datad(alu_io_op2_41),
	.cin(gnd),
	.combout(ShiftRight07),
	.cout());
defparam \ShiftRight0~167 .lut_mask = 16'hAAEE;
defparam \ShiftRight0~167 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~173 (
	.dataa(\_T_60~combout ),
	.datab(\ShiftRight0~172_combout ),
	.datac(gnd),
	.datad(alu_io_op2_41),
	.cin(gnd),
	.combout(ShiftRight08),
	.cout());
defparam \ShiftRight0~173 .lut_mask = 16'hAACC;
defparam \ShiftRight0~173 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~175 (
	.dataa(\ShiftRight0~245_combout ),
	.datab(alu_io_op2_41),
	.datac(\ShiftRight0~174_combout ),
	.datad(\_T_60~combout ),
	.cin(gnd),
	.combout(ShiftRight09),
	.cout());
defparam \ShiftRight0~175 .lut_mask = 16'hF838;
defparam \ShiftRight0~175 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~180 (
	.dataa(\_T_60~combout ),
	.datab(\ShiftRight0~179_combout ),
	.datac(gnd),
	.datad(alu_io_op2_41),
	.cin(gnd),
	.combout(ShiftRight010),
	.cout());
defparam \ShiftRight0~180 .lut_mask = 16'hAACC;
defparam \ShiftRight0~180 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~183 (
	.dataa(\ShiftRight0~243_combout ),
	.datab(alu_io_op2_32),
	.datac(\ShiftRight0~182_combout ),
	.datad(\_T_60~combout ),
	.cin(gnd),
	.combout(ShiftRight011),
	.cout());
defparam \ShiftRight0~183 .lut_mask = 16'hF838;
defparam \ShiftRight0~183 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~188 (
	.dataa(\_T_60~combout ),
	.datab(\ShiftRight0~187_combout ),
	.datac(gnd),
	.datad(alu_io_op2_41),
	.cin(gnd),
	.combout(ShiftRight012),
	.cout());
defparam \ShiftRight0~188 .lut_mask = 16'hAACC;
defparam \ShiftRight0~188 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~190 (
	.dataa(\ShiftRight0~133_combout ),
	.datab(alu_io_op2_41),
	.datac(\ShiftRight0~189_combout ),
	.datad(\_T_60~combout ),
	.cin(gnd),
	.combout(ShiftRight013),
	.cout());
defparam \ShiftRight0~190 .lut_mask = 16'hF838;
defparam \ShiftRight0~190 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~195 (
	.dataa(\_T_60~combout ),
	.datab(\ShiftRight0~194_combout ),
	.datac(gnd),
	.datad(alu_io_op2_41),
	.cin(gnd),
	.combout(ShiftRight014),
	.cout());
defparam \ShiftRight0~195 .lut_mask = 16'hAACC;
defparam \ShiftRight0~195 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~197 (
	.dataa(\ShiftRight0~244_combout ),
	.datab(alu_io_op2_32),
	.datac(\ShiftRight0~196_combout ),
	.datad(\_T_60~combout ),
	.cin(gnd),
	.combout(ShiftRight015),
	.cout());
defparam \ShiftRight0~197 .lut_mask = 16'hF838;
defparam \ShiftRight0~197 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~198 (
	.dataa(\ShiftRight0~248_combout ),
	.datab(alu_io_op2_32),
	.datac(\ShiftRight0~155_combout ),
	.datad(alu_io_op2_41),
	.cin(gnd),
	.combout(ShiftRight016),
	.cout());
defparam \ShiftRight0~198 .lut_mask = 16'hAAEA;
defparam \ShiftRight0~198 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~203 (
	.dataa(\ShiftRight0~241_combout ),
	.datab(\ShiftRight0~199_combout ),
	.datac(\ShiftRight0~202_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(ShiftRight017),
	.cout());
defparam \ShiftRight0~203 .lut_mask = 16'hECEC;
defparam \ShiftRight0~203 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_123[13] (
	.dataa(alu_io_op2_3),
	.datab(ex_reg_rs2_bypass_131),
	.datac(alu_io_op2_13),
	.datad(alu_io_op1_131),
	.cin(gnd),
	.combout(_T_123_13),
	.cout());
defparam \_T_123[13] .lut_mask = 16'h07F8;
defparam \_T_123[13] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~209 (
	.dataa(\ShiftRight0~205_combout ),
	.datab(\ShiftRight0~208_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(ShiftRight018),
	.cout());
defparam \ShiftRight0~209 .lut_mask = 16'hEEEE;
defparam \ShiftRight0~209 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~216 (
	.dataa(\ShiftRight0~241_combout ),
	.datab(\ShiftRight0~212_combout ),
	.datac(\ShiftRight0~215_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(ShiftRight019),
	.cout());
defparam \ShiftRight0~216 .lut_mask = 16'hECEC;
defparam \ShiftRight0~216 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~217 (
	.dataa(alu_io_op2_41),
	.datab(\ShiftRight0~241_combout ),
	.datac(\ShiftRight0~108_combout ),
	.datad(\_T_60~combout ),
	.cin(gnd),
	.combout(ShiftRight020),
	.cout());
defparam \ShiftRight0~217 .lut_mask = 16'hEAC0;
defparam \ShiftRight0~217 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~222 (
	.dataa(\ShiftRight0~218_combout ),
	.datab(\ShiftRight0~221_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(ShiftRight021),
	.cout());
defparam \ShiftRight0~222 .lut_mask = 16'hEEEE;
defparam \ShiftRight0~222 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_139[18] (
	.dataa(alu_io_op1_181),
	.datab(alu_io_op2_18),
	.datac(alu_io_op2_3),
	.datad(ex_reg_rs2_bypass_18),
	.cin(gnd),
	.combout(_T_139_18),
	.cout());
defparam \_T_139[18] .lut_mask = 16'hFEEE;
defparam \_T_139[18] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~228 (
	.dataa(\ShiftRight0~223_combout ),
	.datab(\ShiftRight0~225_combout ),
	.datac(\ShiftRight0~227_combout ),
	.datad(\ShiftRight0~194_combout ),
	.cin(gnd),
	.combout(ShiftRight022),
	.cout());
defparam \ShiftRight0~228 .lut_mask = 16'hF838;
defparam \ShiftRight0~228 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~233 (
	.dataa(\ShiftRight0~229_combout ),
	.datab(\ShiftRight0~37_combout ),
	.datac(\ShiftRight0~232_combout ),
	.datad(\ShiftRight0~187_combout ),
	.cin(gnd),
	.combout(ShiftRight023),
	.cout());
defparam \ShiftRight0~233 .lut_mask = 16'hF2C2;
defparam \ShiftRight0~233 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~236 (
	.dataa(\ShiftRight0~234_combout ),
	.datab(\ShiftRight0~225_combout ),
	.datac(\ShiftRight0~235_combout ),
	.datad(\ShiftRight0~179_combout ),
	.cin(gnd),
	.combout(ShiftRight024),
	.cout());
defparam \ShiftRight0~236 .lut_mask = 16'hF838;
defparam \ShiftRight0~236 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~240 (
	.dataa(\ShiftRight0~237_combout ),
	.datab(\ShiftRight0~37_combout ),
	.datac(\ShiftRight0~239_combout ),
	.datad(\ShiftRight0~172_combout ),
	.cin(gnd),
	.combout(ShiftRight025),
	.cout());
defparam \ShiftRight0~240 .lut_mask = 16'hF2C2;
defparam \ShiftRight0~240 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_123[23] (
	.dataa(ex_ctrl_alu_op1_0),
	.datab(ex_ctrl_alu_op1_1),
	.datac(alu_io_op2_23),
	.datad(alu_io_op1_23),
	.cin(gnd),
	.combout(_T_123_23),
	.cout());
defparam \_T_123[23] .lut_mask = 16'h96F0;
defparam \_T_123[23] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_123[27] (
	.dataa(ex_ctrl_alu_op1_0),
	.datab(ex_ctrl_alu_op1_1),
	.datac(alu_io_op2_27),
	.datad(alu_io_op1_27),
	.cin(gnd),
	.combout(_T_123_27),
	.cout());
defparam \_T_123[27] .lut_mask = 16'h96F0;
defparam \_T_123[27] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_123[29] (
	.dataa(ex_ctrl_alu_op1_0),
	.datab(ex_ctrl_alu_op1_1),
	.datac(alu_io_op2_29),
	.datad(alu_io_op1_29),
	.cin(gnd),
	.combout(_T_123_29),
	.cout());
defparam \_T_123[29] .lut_mask = 16'h96F0;
defparam \_T_123[29] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~249 (
	.dataa(alu_io_op2_32),
	.datab(alu_io_op2_41),
	.datac(\ShiftRight0~204_combout ),
	.datad(\ShiftRight0~139_combout ),
	.cin(gnd),
	.combout(ShiftRight026),
	.cout());
defparam \ShiftRight0~249 .lut_mask = 16'hF1F0;
defparam \ShiftRight0~249 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~250 (
	.dataa(alu_io_op2_32),
	.datab(alu_io_op2_41),
	.datac(\ShiftRight0~210_combout ),
	.datad(\ShiftRight0~243_combout ),
	.cin(gnd),
	.combout(ShiftRight027),
	.cout());
defparam \ShiftRight0~250 .lut_mask = 16'hF1F0;
defparam \ShiftRight0~250 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_123[17] (
	.dataa(ex_ctrl_alu_op1_0),
	.datab(ex_ctrl_alu_op1_1),
	.datac(alu_io_op2_171),
	.datad(alu_io_op1_17),
	.cin(gnd),
	.combout(_T_123_17),
	.cout());
defparam \_T_123[17] .lut_mask = 16'h96F0;
defparam \_T_123[17] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~251 (
	.dataa(alu_io_op2_32),
	.datab(alu_io_op2_41),
	.datac(\ShiftRight0~155_combout ),
	.datad(\_T_60~combout ),
	.cin(gnd),
	.combout(ShiftRight028),
	.cout());
defparam \ShiftRight0~251 .lut_mask = 16'hFE10;
defparam \ShiftRight0~251 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~253 (
	.dataa(alu_io_op2_32),
	.datab(alu_io_op2_41),
	.datac(\ShiftRight0~133_combout ),
	.datad(\_T_60~combout ),
	.cin(gnd),
	.combout(ShiftRight029),
	.cout());
defparam \ShiftRight0~253 .lut_mask = 16'hFE10;
defparam \ShiftRight0~253 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~254 (
	.dataa(alu_io_op2_32),
	.datab(alu_io_op2_41),
	.datac(\ShiftRight0~78_combout ),
	.datad(\_T_60~combout ),
	.cin(gnd),
	.combout(ShiftRight030),
	.cout());
defparam \ShiftRight0~254 .lut_mask = 16'hFE10;
defparam \ShiftRight0~254 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~256 (
	.dataa(alu_io_op2_32),
	.datab(alu_io_op2_41),
	.datac(\ShiftRight0~245_combout ),
	.datad(\_T_60~combout ),
	.cin(gnd),
	.combout(ShiftRight031),
	.cout());
defparam \ShiftRight0~256 .lut_mask = 16'hFE10;
defparam \ShiftRight0~256 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_123[21] (
	.dataa(ex_ctrl_alu_op1_0),
	.datab(ex_ctrl_alu_op1_1),
	.datac(alu_io_op2_21),
	.datad(alu_io_op1_21),
	.cin(gnd),
	.combout(_T_123_21),
	.cout());
defparam \_T_123[21] .lut_mask = 16'h96F0;
defparam \_T_123[21] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_123[25] (
	.dataa(ex_ctrl_alu_op1_0),
	.datab(ex_ctrl_alu_op1_1),
	.datac(alu_io_op2_25),
	.datad(alu_io_op1_25),
	.cin(gnd),
	.combout(_T_123_25),
	.cout());
defparam \_T_123[25] .lut_mask = 16'h96F0;
defparam \_T_123[25] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[0]~46 (
	.dataa(ex_ctrl_alu_op201),
	.datab(ex_ctrl_alu_op210),
	.datac(csr_io_alu_op2_0),
	.datad(ex_reg_rs2_bypass_0),
	.cin(gnd),
	.combout(\op2_inv[0]~46_combout ),
	.cout());
defparam \op2_inv[0]~46 .lut_mask = 16'h070F;
defparam \op2_inv[0]~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[0]~42 (
	.dataa(ex_ctrl_alu_func_3),
	.datab(alu_io_op2_3),
	.datac(ex_reg_rs2_bypass_01),
	.datad(\op2_inv[0]~46_combout ),
	.cin(gnd),
	.combout(\op2_inv[0]~42_combout ),
	.cout());
defparam \op2_inv[0]~42 .lut_mask = 16'h6A55;
defparam \op2_inv[0]~42 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Add0~1 (
	.dataa(ex_ctrl_alu_func_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add0~1_cout ));
defparam \Add0~1 .lut_mask = 16'h00AA;
defparam \Add0~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[1]~45 (
	.dataa(ex_ctrl_alu_op201),
	.datab(ex_ctrl_alu_op210),
	.datac(ex_ctrl_imm_type011),
	.datad(io_sw_r_ex_imm_1),
	.cin(gnd),
	.combout(\op2_inv[1]~45_combout ),
	.cout());
defparam \op2_inv[1]~45 .lut_mask = 16'h7477;
defparam \op2_inv[1]~45 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[1]~41 (
	.dataa(ex_ctrl_alu_func_3),
	.datab(ex_reg_rs2_bypass_1),
	.datac(ex_ctrl_alu_op210),
	.datad(\op2_inv[1]~45_combout ),
	.cin(gnd),
	.combout(\op2_inv[1]~41_combout ),
	.cout());
defparam \op2_inv[1]~41 .lut_mask = 16'hAA65;
defparam \op2_inv[1]~41 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[2]~40 (
	.dataa(gnd),
	.datab(ex_ctrl_alu_func_3),
	.datac(csr_io_alu_op2_1),
	.datad(alu_io_op2_2),
	.cin(gnd),
	.combout(\op2_inv[2]~40_combout ),
	.cout());
defparam \op2_inv[2]~40 .lut_mask = 16'h3CCC;
defparam \op2_inv[2]~40 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[3]~38 (
	.dataa(io_sw_r_ex_imm_3),
	.datab(ex_ctrl_alu_op210),
	.datac(ex_ctrl_imm_type011),
	.datad(gnd),
	.cin(gnd),
	.combout(\op2_inv[3]~38_combout ),
	.cout());
defparam \op2_inv[3]~38 .lut_mask = 16'hFDFD;
defparam \op2_inv[3]~38 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[3]~39 (
	.dataa(ex_ctrl_alu_func_3),
	.datab(alu_io_op2_31),
	.datac(\op2_inv[3]~38_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\op2_inv[3]~39_combout ),
	.cout());
defparam \op2_inv[3]~39 .lut_mask = 16'h6565;
defparam \op2_inv[3]~39 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[4]~36 (
	.dataa(io_sw_r_ex_imm_4),
	.datab(ex_ctrl_alu_op210),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\op2_inv[4]~36_combout ),
	.cout());
defparam \op2_inv[4]~36 .lut_mask = 16'hDDDD;
defparam \op2_inv[4]~36 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[4]~37 (
	.dataa(ex_ctrl_alu_func_3),
	.datab(csr_io_alu_op2_1),
	.datac(alu_io_op2_4),
	.datad(\op2_inv[4]~36_combout ),
	.cin(gnd),
	.combout(\op2_inv[4]~37_combout ),
	.cout());
defparam \op2_inv[4]~37 .lut_mask = 16'h6A66;
defparam \op2_inv[4]~37 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[5]~35 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_5),
	.cin(gnd),
	.combout(\op2_inv[5]~35_combout ),
	.cout());
defparam \op2_inv[5]~35 .lut_mask = 16'h0FF0;
defparam \op2_inv[5]~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[6]~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_6),
	.cin(gnd),
	.combout(\op2_inv[6]~34_combout ),
	.cout());
defparam \op2_inv[6]~34 .lut_mask = 16'h0FF0;
defparam \op2_inv[6]~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[7]~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_7),
	.cin(gnd),
	.combout(\op2_inv[7]~33_combout ),
	.cout());
defparam \op2_inv[7]~33 .lut_mask = 16'h0FF0;
defparam \op2_inv[7]~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[8]~32 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_8),
	.cin(gnd),
	.combout(\op2_inv[8]~32_combout ),
	.cout());
defparam \op2_inv[8]~32 .lut_mask = 16'h0FF0;
defparam \op2_inv[8]~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[9]~31 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_9),
	.cin(gnd),
	.combout(\op2_inv[9]~31_combout ),
	.cout());
defparam \op2_inv[9]~31 .lut_mask = 16'h0FF0;
defparam \op2_inv[9]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[10]~30 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_10),
	.cin(gnd),
	.combout(\op2_inv[10]~30_combout ),
	.cout());
defparam \op2_inv[10]~30 .lut_mask = 16'h0FF0;
defparam \op2_inv[10]~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[11]~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_11),
	.cin(gnd),
	.combout(\op2_inv[11]~29_combout ),
	.cout());
defparam \op2_inv[11]~29 .lut_mask = 16'h0FF0;
defparam \op2_inv[11]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[12]~27 (
	.dataa(alu_io_op2_3),
	.datab(alu_io_op2_12),
	.datac(_T_3681),
	.datad(mem_csr_data_12),
	.cin(gnd),
	.combout(\op2_inv[12]~27_combout ),
	.cout());
defparam \op2_inv[12]~27 .lut_mask = 16'h1333;
defparam \op2_inv[12]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[12]~28 (
	.dataa(alu_io_op2_3),
	.datab(ex_ctrl_alu_func_3),
	.datac(ex_reg_rs2_bypass_12),
	.datad(\op2_inv[12]~27_combout ),
	.cin(gnd),
	.combout(\op2_inv[12]~28_combout ),
	.cout());
defparam \op2_inv[12]~28 .lut_mask = 16'h6C33;
defparam \op2_inv[12]~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[13]~25 (
	.dataa(alu_io_op2_3),
	.datab(alu_io_op2_13),
	.datac(_T_3681),
	.datad(mem_csr_data_13),
	.cin(gnd),
	.combout(\op2_inv[13]~25_combout ),
	.cout());
defparam \op2_inv[13]~25 .lut_mask = 16'h1333;
defparam \op2_inv[13]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[13]~26 (
	.dataa(alu_io_op2_3),
	.datab(ex_ctrl_alu_func_3),
	.datac(ex_reg_rs2_bypass_13),
	.datad(\op2_inv[13]~25_combout ),
	.cin(gnd),
	.combout(\op2_inv[13]~26_combout ),
	.cout());
defparam \op2_inv[13]~26 .lut_mask = 16'h6C33;
defparam \op2_inv[13]~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[14]~23 (
	.dataa(alu_io_op2_3),
	.datab(alu_io_op2_14),
	.datac(_T_3681),
	.datad(mem_csr_data_14),
	.cin(gnd),
	.combout(\op2_inv[14]~23_combout ),
	.cout());
defparam \op2_inv[14]~23 .lut_mask = 16'h1333;
defparam \op2_inv[14]~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[14]~24 (
	.dataa(alu_io_op2_3),
	.datab(ex_ctrl_alu_func_3),
	.datac(ex_reg_rs2_bypass_14),
	.datad(\op2_inv[14]~23_combout ),
	.cin(gnd),
	.combout(\op2_inv[14]~24_combout ),
	.cout());
defparam \op2_inv[14]~24 .lut_mask = 16'h6C33;
defparam \op2_inv[14]~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[15]~22 (
	.dataa(alu_io_op2_3),
	.datab(ex_reg_rs2_bypass_15),
	.datac(alu_io_op2_15),
	.datad(ex_ctrl_alu_func_3),
	.cin(gnd),
	.combout(\op2_inv[15]~22_combout ),
	.cout());
defparam \op2_inv[15]~22 .lut_mask = 16'h07F8;
defparam \op2_inv[15]~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[16]~21 (
	.dataa(alu_io_op2_3),
	.datab(ex_reg_rs2_bypass_16),
	.datac(alu_io_op2_16),
	.datad(ex_ctrl_alu_func_3),
	.cin(gnd),
	.combout(\op2_inv[16]~21_combout ),
	.cout());
defparam \op2_inv[16]~21 .lut_mask = 16'h07F8;
defparam \op2_inv[16]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[17]~20 (
	.dataa(alu_io_op2_3),
	.datab(ex_reg_rs2_bypass_17),
	.datac(alu_io_op2_17),
	.datad(ex_ctrl_alu_func_3),
	.cin(gnd),
	.combout(\op2_inv[17]~20_combout ),
	.cout());
defparam \op2_inv[17]~20 .lut_mask = 16'h07F8;
defparam \op2_inv[17]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[18]~19 (
	.dataa(alu_io_op2_3),
	.datab(ex_reg_rs2_bypass_18),
	.datac(alu_io_op2_18),
	.datad(ex_ctrl_alu_func_3),
	.cin(gnd),
	.combout(\op2_inv[18]~19_combout ),
	.cout());
defparam \op2_inv[18]~19 .lut_mask = 16'h07F8;
defparam \op2_inv[18]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[19]~18 (
	.dataa(alu_io_op2_3),
	.datab(ex_reg_rs2_bypass_19),
	.datac(alu_io_op2_19),
	.datad(ex_ctrl_alu_func_3),
	.cin(gnd),
	.combout(\op2_inv[19]~18_combout ),
	.cout());
defparam \op2_inv[19]~18 .lut_mask = 16'h07F8;
defparam \op2_inv[19]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[20]~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_20),
	.cin(gnd),
	.combout(\op2_inv[20]~17_combout ),
	.cout());
defparam \op2_inv[20]~17 .lut_mask = 16'h0FF0;
defparam \op2_inv[20]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[21]~16 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_21),
	.cin(gnd),
	.combout(\op2_inv[21]~16_combout ),
	.cout());
defparam \op2_inv[21]~16 .lut_mask = 16'h0FF0;
defparam \op2_inv[21]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[22]~15 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_22),
	.cin(gnd),
	.combout(\op2_inv[22]~15_combout ),
	.cout());
defparam \op2_inv[22]~15 .lut_mask = 16'h0FF0;
defparam \op2_inv[22]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[23]~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_23),
	.cin(gnd),
	.combout(\op2_inv[23]~14_combout ),
	.cout());
defparam \op2_inv[23]~14 .lut_mask = 16'h0FF0;
defparam \op2_inv[23]~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[24]~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_24),
	.cin(gnd),
	.combout(\op2_inv[24]~13_combout ),
	.cout());
defparam \op2_inv[24]~13 .lut_mask = 16'h0FF0;
defparam \op2_inv[24]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[25]~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_25),
	.cin(gnd),
	.combout(\op2_inv[25]~12_combout ),
	.cout());
defparam \op2_inv[25]~12 .lut_mask = 16'h0FF0;
defparam \op2_inv[25]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[26]~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_26),
	.cin(gnd),
	.combout(\op2_inv[26]~11_combout ),
	.cout());
defparam \op2_inv[26]~11 .lut_mask = 16'h0FF0;
defparam \op2_inv[26]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[27]~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_27),
	.cin(gnd),
	.combout(\op2_inv[27]~10_combout ),
	.cout());
defparam \op2_inv[27]~10 .lut_mask = 16'h0FF0;
defparam \op2_inv[27]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[28]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_28),
	.cin(gnd),
	.combout(\op2_inv[28]~9_combout ),
	.cout());
defparam \op2_inv[28]~9 .lut_mask = 16'h0FF0;
defparam \op2_inv[28]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[29]~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_29),
	.cin(gnd),
	.combout(\op2_inv[29]~8_combout ),
	.cout());
defparam \op2_inv[29]~8 .lut_mask = 16'h0FF0;
defparam \op2_inv[29]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[30]~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_30),
	.cin(gnd),
	.combout(\op2_inv[30]~7_combout ),
	.cout());
defparam \op2_inv[30]~7 .lut_mask = 16'h0FF0;
defparam \op2_inv[30]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[31]~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ex_ctrl_alu_func_3),
	.datad(alu_io_op2_311),
	.cin(gnd),
	.combout(\op2_inv[31]~6_combout ),
	.cout());
defparam \op2_inv[31]~6 .lut_mask = 16'h0FF0;
defparam \op2_inv[31]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~0 (
	.dataa(alu_io_op1_281),
	.datab(alu_io_op1_291),
	.datac(alu_io_op2_29),
	.datad(alu_io_op2_28),
	.cin(gnd),
	.combout(\_T_125~0_combout ),
	.cout());
defparam \_T_125~0 .lut_mask = 16'h8241;
defparam \_T_125~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~1 (
	.dataa(\_T_125~0_combout ),
	.datab(alu_io_op1_301),
	.datac(alu_io_op2_30),
	.datad(_T_123_31),
	.cin(gnd),
	.combout(\_T_125~1_combout ),
	.cout());
defparam \_T_125~1 .lut_mask = 16'h0082;
defparam \_T_125~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~2 (
	.dataa(csr_io_alu_op2_01),
	.datab(csr_io_alu_op1_11),
	.datac(csr_io_alu_op2_11),
	.datad(csr_io_alu_op1_02),
	.cin(gnd),
	.combout(\_T_125~2_combout ),
	.cout());
defparam \_T_125~2 .lut_mask = 16'h8241;
defparam \_T_125~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~3 (
	.dataa(alu_io_op1_81),
	.datab(alu_io_op1_91),
	.datac(alu_io_op2_9),
	.datad(alu_io_op2_8),
	.cin(gnd),
	.combout(\_T_125~3_combout ),
	.cout());
defparam \_T_125~3 .lut_mask = 16'h8241;
defparam \_T_125~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~4 (
	.dataa(\_T_125~3_combout ),
	.datab(alu_io_op1_101),
	.datac(alu_io_op2_10),
	.datad(_T_123_11),
	.cin(gnd),
	.combout(\_T_125~4_combout ),
	.cout());
defparam \_T_125~4 .lut_mask = 16'h0082;
defparam \_T_125~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~5 (
	.dataa(alu_io_op1_121),
	.datab(alu_io_op1_131),
	.datac(alu_io_op2_131),
	.datad(alu_io_op2_121),
	.cin(gnd),
	.combout(\_T_125~5_combout ),
	.cout());
defparam \_T_125~5 .lut_mask = 16'h8241;
defparam \_T_125~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~6 (
	.dataa(\_T_125~5_combout ),
	.datab(alu_io_op1_141),
	.datac(alu_io_op2_141),
	.datad(_T_123_15),
	.cin(gnd),
	.combout(\_T_125~6_combout ),
	.cout());
defparam \_T_125~6 .lut_mask = 16'h0082;
defparam \_T_125~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~7 (
	.dataa(alu_io_op1_161),
	.datab(alu_io_op1_171),
	.datac(alu_io_op2_171),
	.datad(alu_io_op2_161),
	.cin(gnd),
	.combout(\_T_125~7_combout ),
	.cout());
defparam \_T_125~7 .lut_mask = 16'h8241;
defparam \_T_125~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~8 (
	.dataa(\_T_125~7_combout ),
	.datab(alu_io_op1_181),
	.datac(alu_io_op2_181),
	.datad(_T_123_19),
	.cin(gnd),
	.combout(\_T_125~8_combout ),
	.cout());
defparam \_T_125~8 .lut_mask = 16'h0082;
defparam \_T_125~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~9 (
	.dataa(\_T_125~2_combout ),
	.datab(\_T_125~4_combout ),
	.datac(\_T_125~6_combout ),
	.datad(\_T_125~8_combout ),
	.cin(gnd),
	.combout(\_T_125~9_combout ),
	.cout());
defparam \_T_125~9 .lut_mask = 16'h8000;
defparam \_T_125~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~10 (
	.dataa(alu_io_op2_41),
	.datab(alu_io_op1_41),
	.datac(ex_ctrl_alu_func_3),
	.datad(_T_123_2),
	.cin(gnd),
	.combout(\_T_125~10_combout ),
	.cout());
defparam \_T_125~10 .lut_mask = 16'h0009;
defparam \_T_125~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~11 (
	.dataa(alu_io_op2_32),
	.datab(alu_io_op1_51),
	.datac(alu_io_op2_5),
	.datad(alu_io_op1_32),
	.cin(gnd),
	.combout(\_T_125~11_combout ),
	.cout());
defparam \_T_125~11 .lut_mask = 16'h8241;
defparam \_T_125~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~12 (
	.dataa(\_T_125~11_combout ),
	.datab(alu_io_op1_61),
	.datac(alu_io_op2_6),
	.datad(_T_123_7),
	.cin(gnd),
	.combout(\_T_125~12_combout ),
	.cout());
defparam \_T_125~12 .lut_mask = 16'h0082;
defparam \_T_125~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~13 (
	.dataa(alu_io_op1_201),
	.datab(alu_io_op1_211),
	.datac(alu_io_op2_21),
	.datad(alu_io_op2_20),
	.cin(gnd),
	.combout(\_T_125~13_combout ),
	.cout());
defparam \_T_125~13 .lut_mask = 16'h8241;
defparam \_T_125~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~14 (
	.dataa(\_T_125~13_combout ),
	.datab(alu_io_op1_221),
	.datac(alu_io_op2_22),
	.datad(_T_123_23),
	.cin(gnd),
	.combout(\_T_125~14_combout ),
	.cout());
defparam \_T_125~14 .lut_mask = 16'h0082;
defparam \_T_125~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~15 (
	.dataa(alu_io_op1_241),
	.datab(alu_io_op1_251),
	.datac(alu_io_op2_25),
	.datad(alu_io_op2_24),
	.cin(gnd),
	.combout(\_T_125~15_combout ),
	.cout());
defparam \_T_125~15 .lut_mask = 16'h8241;
defparam \_T_125~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~16 (
	.dataa(\_T_125~15_combout ),
	.datab(alu_io_op1_261),
	.datac(alu_io_op2_26),
	.datad(_T_123_27),
	.cin(gnd),
	.combout(\_T_125~16_combout ),
	.cout());
defparam \_T_125~16 .lut_mask = 16'h0082;
defparam \_T_125~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~17 (
	.dataa(\_T_125~10_combout ),
	.datab(\_T_125~12_combout ),
	.datac(\_T_125~14_combout ),
	.datad(\_T_125~16_combout ),
	.cin(gnd),
	.combout(\_T_125~17_combout ),
	.cout());
defparam \_T_125~17 .lut_mask = 16'h8000;
defparam \_T_125~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~18 (
	.dataa(ex_ctrl_alu_func_3),
	.datab(alu_io_op1_311),
	.datac(LessThan0),
	.datad(alu_io_op2_311),
	.cin(gnd),
	.combout(\_T_125~18_combout ),
	.cout());
defparam \_T_125~18 .lut_mask = 16'h0280;
defparam \_T_125~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_125~19 (
	.dataa(ex_ctrl_alu_func_3),
	.datab(_T_123_31),
	.datac(\_T_125~18_combout ),
	.datad(_T_3_31),
	.cin(gnd),
	.combout(\_T_125~19_combout ),
	.cout());
defparam \_T_125~19 .lut_mask = 16'hF2F0;
defparam \_T_125~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~241 (
	.dataa(ex_ctrl_alu_op1_0),
	.datab(ex_ctrl_alu_op1_1),
	.datac(alu_io_op2_41),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~241_combout ),
	.cout());
defparam \ShiftRight0~241 .lut_mask = 16'h0606;
defparam \ShiftRight0~241 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_8~0 (
	.dataa(ex_ctrl_alu_func_3),
	.datab(ex_ctrl_alu_func_2),
	.datac(ex_ctrl_alu_func_1),
	.datad(ex_ctrl_alu_func_0),
	.cin(gnd),
	.combout(\_T_8~0_combout ),
	.cout());
defparam \_T_8~0 .lut_mask = 16'h2400;
defparam \_T_8~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~32 (
	.dataa(csr_io_alu_op2_01),
	.datab(alu_io_op1_31),
	.datac(csr_io_alu_op1_01),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~32_combout ),
	.cout());
defparam \ShiftRight0~32 .lut_mask = 16'h88A0;
defparam \ShiftRight0~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~33 (
	.dataa(alu_io_op1_30),
	.datab(csr_io_alu_op1_1),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~33_combout ),
	.cout());
defparam \ShiftRight0~33 .lut_mask = 16'hAACC;
defparam \ShiftRight0~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~34 (
	.dataa(\ShiftRight0~32_combout ),
	.datab(\ShiftRight0~33_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~34_combout ),
	.cout());
defparam \ShiftRight0~34 .lut_mask = 16'hAAEE;
defparam \ShiftRight0~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~35 (
	.dataa(alu_io_op2_2),
	.datab(ex_reg_rs2_bypass_1),
	.datac(io_sw_r_ex_imm_1),
	.datad(ex_ctrl_alu_op210),
	.cin(gnd),
	.combout(\ShiftRight0~35_combout ),
	.cout());
defparam \ShiftRight0~35 .lut_mask = 16'hEEFA;
defparam \ShiftRight0~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~242 (
	.dataa(ex_ctrl_alu_op201),
	.datab(ex_ctrl_alu_op210),
	.datac(ex_ctrl_imm_type011),
	.datad(\ShiftRight0~35_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~242_combout ),
	.cout());
defparam \ShiftRight0~242 .lut_mask = 16'h8B00;
defparam \ShiftRight0~242 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~36 (
	.dataa(\ShiftRight0~241_combout ),
	.datab(\ShiftRight0~34_combout ),
	.datac(alu_io_op2_32),
	.datad(\ShiftRight0~242_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~36_combout ),
	.cout());
defparam \ShiftRight0~36 .lut_mask = 16'h0008;
defparam \ShiftRight0~36 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb _T_60(
	.dataa(ex_ctrl_alu_func_3),
	.datab(alu_io_op1_311),
	.datac(csr_io_alu_op1_02),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\_T_60~combout ),
	.cout());
defparam _T_60.lut_mask = 16'h88A0;
defparam _T_60.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(alu_io_op2_32),
	.datad(alu_io_op2_41),
	.cin(gnd),
	.combout(\ShiftRight0~37_combout ),
	.cout());
defparam \ShiftRight0~37 .lut_mask = 16'h000F;
defparam \ShiftRight0~37 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~39 (
	.dataa(alu_io_op1_8),
	.datab(alu_io_op1_23),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~39_combout ),
	.cout());
defparam \ShiftRight0~39 .lut_mask = 16'hAACC;
defparam \ShiftRight0~39 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~40 (
	.dataa(alu_io_op1_7),
	.datab(alu_io_op1_24),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~40_combout ),
	.cout());
defparam \ShiftRight0~40 .lut_mask = 16'hAACC;
defparam \ShiftRight0~40 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~41 (
	.dataa(\ShiftRight0~39_combout ),
	.datab(\ShiftRight0~40_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~41_combout ),
	.cout());
defparam \ShiftRight0~41 .lut_mask = 16'hAACC;
defparam \ShiftRight0~41 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~42 (
	.dataa(alu_io_op1_4),
	.datab(alu_io_op1_27),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~42_combout ),
	.cout());
defparam \ShiftRight0~42 .lut_mask = 16'hAACC;
defparam \ShiftRight0~42 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~43 (
	.dataa(alu_io_op1_3),
	.datab(alu_io_op1_28),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~43_combout ),
	.cout());
defparam \ShiftRight0~43 .lut_mask = 16'hAACC;
defparam \ShiftRight0~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~44 (
	.dataa(\ShiftRight0~42_combout ),
	.datab(\ShiftRight0~43_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~44_combout ),
	.cout());
defparam \ShiftRight0~44 .lut_mask = 16'hAACC;
defparam \ShiftRight0~44 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~45 (
	.dataa(csr_io_alu_op2_11),
	.datab(\ShiftRight0~41_combout ),
	.datac(\ShiftRight0~44_combout ),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~45_combout ),
	.cout());
defparam \ShiftRight0~45 .lut_mask = 16'h88A0;
defparam \ShiftRight0~45 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~46 (
	.dataa(alu_io_op1_6),
	.datab(alu_io_op1_25),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~46_combout ),
	.cout());
defparam \ShiftRight0~46 .lut_mask = 16'hAACC;
defparam \ShiftRight0~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~47 (
	.dataa(alu_io_op1_5),
	.datab(alu_io_op1_26),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~47_combout ),
	.cout());
defparam \ShiftRight0~47 .lut_mask = 16'hAACC;
defparam \ShiftRight0~47 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~48 (
	.dataa(\ShiftRight0~46_combout ),
	.datab(\ShiftRight0~47_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~48_combout ),
	.cout());
defparam \ShiftRight0~48 .lut_mask = 16'hAACC;
defparam \ShiftRight0~48 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~49 (
	.dataa(\_T_8~0_combout ),
	.datab(alu_io_op1_2),
	.datac(csr_io_alu_op1_1),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~49_combout ),
	.cout());
defparam \ShiftRight0~49 .lut_mask = 16'h88A0;
defparam \ShiftRight0~49 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~50 (
	.dataa(alu_io_op1_29),
	.datab(alu_io_op1_30),
	.datac(csr_io_alu_op2_01),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~50_combout ),
	.cout());
defparam \ShiftRight0~50 .lut_mask = 16'h00AC;
defparam \ShiftRight0~50 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~51 (
	.dataa(\ShiftRight0~48_combout ),
	.datab(\ShiftRight0~49_combout ),
	.datac(\ShiftRight0~50_combout ),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~51_combout ),
	.cout());
defparam \ShiftRight0~51 .lut_mask = 16'hAAFC;
defparam \ShiftRight0~51 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~52 (
	.dataa(\ShiftRight0~45_combout ),
	.datab(\ShiftRight0~51_combout ),
	.datac(csr_io_alu_op2_11),
	.datad(alu_io_op2_32),
	.cin(gnd),
	.combout(\ShiftRight0~52_combout ),
	.cout());
defparam \ShiftRight0~52 .lut_mask = 16'h00AE;
defparam \ShiftRight0~52 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~53 (
	.dataa(alu_io_op1_12),
	.datab(alu_io_op1_19),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~53_combout ),
	.cout());
defparam \ShiftRight0~53 .lut_mask = 16'hAACC;
defparam \ShiftRight0~53 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~54 (
	.dataa(alu_io_op1_11),
	.datab(alu_io_op1_20),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~54_combout ),
	.cout());
defparam \ShiftRight0~54 .lut_mask = 16'hAACC;
defparam \ShiftRight0~54 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~55 (
	.dataa(\ShiftRight0~53_combout ),
	.datab(\ShiftRight0~54_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~55_combout ),
	.cout());
defparam \ShiftRight0~55 .lut_mask = 16'hAACC;
defparam \ShiftRight0~55 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~56 (
	.dataa(alu_io_op1_10),
	.datab(alu_io_op1_21),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~56_combout ),
	.cout());
defparam \ShiftRight0~56 .lut_mask = 16'hAACC;
defparam \ShiftRight0~56 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~57 (
	.dataa(alu_io_op1_9),
	.datab(alu_io_op1_22),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~57_combout ),
	.cout());
defparam \ShiftRight0~57 .lut_mask = 16'hAACC;
defparam \ShiftRight0~57 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~58 (
	.dataa(\ShiftRight0~56_combout ),
	.datab(\ShiftRight0~57_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~58_combout ),
	.cout());
defparam \ShiftRight0~58 .lut_mask = 16'hAACC;
defparam \ShiftRight0~58 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~59 (
	.dataa(\ShiftRight0~55_combout ),
	.datab(\ShiftRight0~58_combout ),
	.datac(csr_io_alu_op2_11),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~59_combout ),
	.cout());
defparam \ShiftRight0~59 .lut_mask = 16'h00AC;
defparam \ShiftRight0~59 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~60 (
	.dataa(alu_io_op1_16),
	.datab(alu_io_op1_15),
	.datac(csr_io_alu_op2_01),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~60_combout ),
	.cout());
defparam \ShiftRight0~60 .lut_mask = 16'hACCA;
defparam \ShiftRight0~60 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~61 (
	.dataa(alu_io_op1_14),
	.datab(alu_io_op1_17),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~61_combout ),
	.cout());
defparam \ShiftRight0~61 .lut_mask = 16'hAACC;
defparam \ShiftRight0~61 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~62 (
	.dataa(alu_io_op1_13),
	.datab(alu_io_op1_18),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~62_combout ),
	.cout());
defparam \ShiftRight0~62 .lut_mask = 16'hAACC;
defparam \ShiftRight0~62 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~63 (
	.dataa(\ShiftRight0~61_combout ),
	.datab(\ShiftRight0~62_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~63_combout ),
	.cout());
defparam \ShiftRight0~63 .lut_mask = 16'hAACC;
defparam \ShiftRight0~63 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~64 (
	.dataa(\ShiftRight0~60_combout ),
	.datab(\ShiftRight0~63_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~64_combout ),
	.cout());
defparam \ShiftRight0~64 .lut_mask = 16'hAACC;
defparam \ShiftRight0~64 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~65 (
	.dataa(\ShiftRight0~59_combout ),
	.datab(alu_io_op2_210),
	.datac(\ShiftRight0~64_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~65_combout ),
	.cout());
defparam \ShiftRight0~65 .lut_mask = 16'hEAEA;
defparam \ShiftRight0~65 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~66 (
	.dataa(\ShiftRight0~241_combout ),
	.datab(\ShiftRight0~52_combout ),
	.datac(alu_io_op2_32),
	.datad(\ShiftRight0~65_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~66_combout ),
	.cout());
defparam \ShiftRight0~66 .lut_mask = 16'hA888;
defparam \ShiftRight0~66 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_62[31]~0 (
	.dataa(csr_io_alu_op1_0),
	.datab(alu_io_op1_31),
	.datac(csr_io_alu_op1_01),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\_T_62[31]~0_combout ),
	.cout());
defparam \_T_62[31]~0 .lut_mask = 16'h88A0;
defparam \_T_62[31]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~67 (
	.dataa(csr_io_alu_op2_11),
	.datab(\_T_62[31]~0_combout ),
	.datac(ex_ctrl_alu_func_3),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~67_combout ),
	.cout());
defparam \ShiftRight0~67 .lut_mask = 16'h8088;
defparam \ShiftRight0~67 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~68 (
	.dataa(alu_io_op1_29),
	.datab(alu_io_op1_2),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~68_combout ),
	.cout());
defparam \ShiftRight0~68 .lut_mask = 16'hAACC;
defparam \ShiftRight0~68 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~69 (
	.dataa(\ShiftRight0~33_combout ),
	.datab(\ShiftRight0~68_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~69_combout ),
	.cout());
defparam \ShiftRight0~69 .lut_mask = 16'hAACC;
defparam \ShiftRight0~69 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~70 (
	.dataa(\ShiftRight0~67_combout ),
	.datab(csr_io_alu_op1_0),
	.datac(\ShiftRight0~69_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~70_combout ),
	.cout());
defparam \ShiftRight0~70 .lut_mask = 16'hAAEA;
defparam \ShiftRight0~70 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~71 (
	.dataa(alu_io_op1_28),
	.datab(alu_io_op1_3),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~71_combout ),
	.cout());
defparam \ShiftRight0~71 .lut_mask = 16'hAACC;
defparam \ShiftRight0~71 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~72 (
	.dataa(alu_io_op1_27),
	.datab(alu_io_op1_4),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~72_combout ),
	.cout());
defparam \ShiftRight0~72 .lut_mask = 16'hAACC;
defparam \ShiftRight0~72 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~73 (
	.dataa(\ShiftRight0~71_combout ),
	.datab(\ShiftRight0~72_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~73_combout ),
	.cout());
defparam \ShiftRight0~73 .lut_mask = 16'hAACC;
defparam \ShiftRight0~73 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~74 (
	.dataa(alu_io_op1_26),
	.datab(alu_io_op1_5),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~74_combout ),
	.cout());
defparam \ShiftRight0~74 .lut_mask = 16'hAACC;
defparam \ShiftRight0~74 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~75 (
	.dataa(alu_io_op1_25),
	.datab(alu_io_op1_6),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~75_combout ),
	.cout());
defparam \ShiftRight0~75 .lut_mask = 16'hAACC;
defparam \ShiftRight0~75 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~76 (
	.dataa(\ShiftRight0~74_combout ),
	.datab(\ShiftRight0~75_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~76_combout ),
	.cout());
defparam \ShiftRight0~76 .lut_mask = 16'hAACC;
defparam \ShiftRight0~76 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~77 (
	.dataa(\ShiftRight0~73_combout ),
	.datab(\ShiftRight0~76_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~77_combout ),
	.cout());
defparam \ShiftRight0~77 .lut_mask = 16'hAACC;
defparam \ShiftRight0~77 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~78 (
	.dataa(\ShiftRight0~70_combout ),
	.datab(csr_io_alu_op1_0),
	.datac(\ShiftRight0~77_combout ),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~78_combout ),
	.cout());
defparam \ShiftRight0~78 .lut_mask = 16'hAAC0;
defparam \ShiftRight0~78 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~79 (
	.dataa(alu_io_op1_20),
	.datab(alu_io_op1_11),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~79_combout ),
	.cout());
defparam \ShiftRight0~79 .lut_mask = 16'hAACC;
defparam \ShiftRight0~79 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~80 (
	.dataa(alu_io_op1_19),
	.datab(alu_io_op1_12),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~80_combout ),
	.cout());
defparam \ShiftRight0~80 .lut_mask = 16'hAACC;
defparam \ShiftRight0~80 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~81 (
	.dataa(\ShiftRight0~79_combout ),
	.datab(\ShiftRight0~80_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~81_combout ),
	.cout());
defparam \ShiftRight0~81 .lut_mask = 16'hAACC;
defparam \ShiftRight0~81 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~82 (
	.dataa(alu_io_op1_18),
	.datab(alu_io_op1_13),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~82_combout ),
	.cout());
defparam \ShiftRight0~82 .lut_mask = 16'hAACC;
defparam \ShiftRight0~82 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~83 (
	.dataa(alu_io_op1_17),
	.datab(alu_io_op1_14),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~83_combout ),
	.cout());
defparam \ShiftRight0~83 .lut_mask = 16'hAACC;
defparam \ShiftRight0~83 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~84 (
	.dataa(\ShiftRight0~82_combout ),
	.datab(\ShiftRight0~83_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~84_combout ),
	.cout());
defparam \ShiftRight0~84 .lut_mask = 16'hAACC;
defparam \ShiftRight0~84 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~85 (
	.dataa(\ShiftRight0~81_combout ),
	.datab(\ShiftRight0~84_combout ),
	.datac(csr_io_alu_op2_11),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~85_combout ),
	.cout());
defparam \ShiftRight0~85 .lut_mask = 16'h00AC;
defparam \ShiftRight0~85 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~86 (
	.dataa(alu_io_op1_24),
	.datab(alu_io_op1_7),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~86_combout ),
	.cout());
defparam \ShiftRight0~86 .lut_mask = 16'hAACC;
defparam \ShiftRight0~86 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~87 (
	.dataa(alu_io_op1_23),
	.datab(alu_io_op1_8),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~87_combout ),
	.cout());
defparam \ShiftRight0~87 .lut_mask = 16'hAACC;
defparam \ShiftRight0~87 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~88 (
	.dataa(\ShiftRight0~86_combout ),
	.datab(\ShiftRight0~87_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~88_combout ),
	.cout());
defparam \ShiftRight0~88 .lut_mask = 16'hAACC;
defparam \ShiftRight0~88 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~89 (
	.dataa(alu_io_op1_22),
	.datab(alu_io_op1_9),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~89_combout ),
	.cout());
defparam \ShiftRight0~89 .lut_mask = 16'hAACC;
defparam \ShiftRight0~89 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~90 (
	.dataa(alu_io_op1_21),
	.datab(alu_io_op1_10),
	.datac(gnd),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~90_combout ),
	.cout());
defparam \ShiftRight0~90 .lut_mask = 16'hAACC;
defparam \ShiftRight0~90 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~91 (
	.dataa(\ShiftRight0~89_combout ),
	.datab(\ShiftRight0~90_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~91_combout ),
	.cout());
defparam \ShiftRight0~91 .lut_mask = 16'hAACC;
defparam \ShiftRight0~91 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~92 (
	.dataa(alu_io_op2_210),
	.datab(\ShiftRight0~88_combout ),
	.datac(\ShiftRight0~91_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~92_combout ),
	.cout());
defparam \ShiftRight0~92 .lut_mask = 16'h88A0;
defparam \ShiftRight0~92 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~243 (
	.dataa(ex_ctrl_alu_op1_0),
	.datab(ex_ctrl_alu_op1_1),
	.datac(\ShiftRight0~85_combout ),
	.datad(\ShiftRight0~92_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~243_combout ),
	.cout());
defparam \ShiftRight0~243 .lut_mask = 16'h6660;
defparam \ShiftRight0~243 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~93 (
	.dataa(alu_io_op2_41),
	.datab(\ShiftRight0~78_combout ),
	.datac(\ShiftRight0~243_combout ),
	.datad(alu_io_op2_32),
	.cin(gnd),
	.combout(\ShiftRight0~93_combout ),
	.cout());
defparam \ShiftRight0~93 .lut_mask = 16'h88A0;
defparam \ShiftRight0~93 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~95 (
	.dataa(\ShiftRight0~80_combout ),
	.datab(\ShiftRight0~82_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~95_combout ),
	.cout());
defparam \ShiftRight0~95 .lut_mask = 16'hAACC;
defparam \ShiftRight0~95 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~96 (
	.dataa(alu_io_op1_16),
	.datab(alu_io_op1_15),
	.datac(\_T_8~0_combout ),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~96_combout ),
	.cout());
defparam \ShiftRight0~96 .lut_mask = 16'h00AC;
defparam \ShiftRight0~96 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~97 (
	.dataa(\ShiftRight0~96_combout ),
	.datab(csr_io_alu_op2_01),
	.datac(\ShiftRight0~83_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~97_combout ),
	.cout());
defparam \ShiftRight0~97 .lut_mask = 16'hEAEA;
defparam \ShiftRight0~97 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~98 (
	.dataa(\ShiftRight0~95_combout ),
	.datab(\ShiftRight0~97_combout ),
	.datac(csr_io_alu_op2_11),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~98_combout ),
	.cout());
defparam \ShiftRight0~98 .lut_mask = 16'h00AC;
defparam \ShiftRight0~98 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~99 (
	.dataa(\ShiftRight0~87_combout ),
	.datab(\ShiftRight0~89_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~99_combout ),
	.cout());
defparam \ShiftRight0~99 .lut_mask = 16'hAACC;
defparam \ShiftRight0~99 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~100 (
	.dataa(\ShiftRight0~90_combout ),
	.datab(\ShiftRight0~79_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~100_combout ),
	.cout());
defparam \ShiftRight0~100 .lut_mask = 16'hAACC;
defparam \ShiftRight0~100 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~101 (
	.dataa(alu_io_op2_210),
	.datab(\ShiftRight0~99_combout ),
	.datac(\ShiftRight0~100_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~101_combout ),
	.cout());
defparam \ShiftRight0~101 .lut_mask = 16'h88A0;
defparam \ShiftRight0~101 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~102 (
	.dataa(\ShiftRight0~98_combout ),
	.datab(\ShiftRight0~101_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~102_combout ),
	.cout());
defparam \ShiftRight0~102 .lut_mask = 16'hEEEE;
defparam \ShiftRight0~102 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~103 (
	.dataa(\ShiftRight0~72_combout ),
	.datab(\ShiftRight0~74_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~103_combout ),
	.cout());
defparam \ShiftRight0~103 .lut_mask = 16'hAACC;
defparam \ShiftRight0~103 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~104 (
	.dataa(\ShiftRight0~75_combout ),
	.datab(\ShiftRight0~86_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~104_combout ),
	.cout());
defparam \ShiftRight0~104 .lut_mask = 16'hAACC;
defparam \ShiftRight0~104 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~105 (
	.dataa(\ShiftRight0~103_combout ),
	.datab(\ShiftRight0~104_combout ),
	.datac(csr_io_alu_op2_11),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~105_combout ),
	.cout());
defparam \ShiftRight0~105 .lut_mask = 16'h00AC;
defparam \ShiftRight0~105 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~106 (
	.dataa(\ShiftRight0~68_combout ),
	.datab(\ShiftRight0~71_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~106_combout ),
	.cout());
defparam \ShiftRight0~106 .lut_mask = 16'hAACC;
defparam \ShiftRight0~106 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~107 (
	.dataa(alu_io_op2_210),
	.datab(\ShiftRight0~34_combout ),
	.datac(\ShiftRight0~106_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~107_combout ),
	.cout());
defparam \ShiftRight0~107 .lut_mask = 16'h88A0;
defparam \ShiftRight0~107 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~108 (
	.dataa(\ShiftRight0~102_combout ),
	.datab(alu_io_op2_32),
	.datac(\ShiftRight0~105_combout ),
	.datad(\ShiftRight0~107_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~108_combout ),
	.cout());
defparam \ShiftRight0~108 .lut_mask = 16'hEEE2;
defparam \ShiftRight0~108 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~109 (
	.dataa(\ShiftRight0~54_combout ),
	.datab(\ShiftRight0~56_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~109_combout ),
	.cout());
defparam \ShiftRight0~109 .lut_mask = 16'hAACC;
defparam \ShiftRight0~109 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~110 (
	.dataa(\ShiftRight0~57_combout ),
	.datab(\ShiftRight0~39_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~110_combout ),
	.cout());
defparam \ShiftRight0~110 .lut_mask = 16'hAACC;
defparam \ShiftRight0~110 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~111 (
	.dataa(\ShiftRight0~109_combout ),
	.datab(\ShiftRight0~110_combout ),
	.datac(csr_io_alu_op2_11),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~111_combout ),
	.cout());
defparam \ShiftRight0~111 .lut_mask = 16'h00AC;
defparam \ShiftRight0~111 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~112 (
	.dataa(csr_io_alu_op2_01),
	.datab(alu_io_op1_15),
	.datac(alu_io_op1_16),
	.datad(\_T_8~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~112_combout ),
	.cout());
defparam \ShiftRight0~112 .lut_mask = 16'h88A0;
defparam \ShiftRight0~112 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~113 (
	.dataa(\ShiftRight0~112_combout ),
	.datab(\ShiftRight0~61_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~113_combout ),
	.cout());
defparam \ShiftRight0~113 .lut_mask = 16'hAAEE;
defparam \ShiftRight0~113 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~114 (
	.dataa(\ShiftRight0~62_combout ),
	.datab(\ShiftRight0~53_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~114_combout ),
	.cout());
defparam \ShiftRight0~114 .lut_mask = 16'hAACC;
defparam \ShiftRight0~114 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~115 (
	.dataa(alu_io_op2_210),
	.datab(\ShiftRight0~113_combout ),
	.datac(\ShiftRight0~114_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~115_combout ),
	.cout());
defparam \ShiftRight0~115 .lut_mask = 16'h88A0;
defparam \ShiftRight0~115 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~116 (
	.dataa(\ShiftRight0~111_combout ),
	.datab(\ShiftRight0~115_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~116_combout ),
	.cout());
defparam \ShiftRight0~116 .lut_mask = 16'hEEEE;
defparam \ShiftRight0~116 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~117 (
	.dataa(\ShiftRight0~40_combout ),
	.datab(\ShiftRight0~46_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~117_combout ),
	.cout());
defparam \ShiftRight0~117 .lut_mask = 16'hAACC;
defparam \ShiftRight0~117 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~118 (
	.dataa(alu_io_op1_2),
	.datab(alu_io_op1_29),
	.datac(\_T_8~0_combout ),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~118_combout ),
	.cout());
defparam \ShiftRight0~118 .lut_mask = 16'h00AC;
defparam \ShiftRight0~118 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~119 (
	.dataa(\ShiftRight0~118_combout ),
	.datab(csr_io_alu_op2_01),
	.datac(\ShiftRight0~43_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~119_combout ),
	.cout());
defparam \ShiftRight0~119 .lut_mask = 16'hEAEA;
defparam \ShiftRight0~119 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~120 (
	.dataa(csr_io_alu_op2_11),
	.datab(\ShiftRight0~117_combout ),
	.datac(\ShiftRight0~119_combout ),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~120_combout ),
	.cout());
defparam \ShiftRight0~120 .lut_mask = 16'h88A0;
defparam \ShiftRight0~120 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~121 (
	.dataa(\ShiftRight0~47_combout ),
	.datab(\ShiftRight0~42_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~121_combout ),
	.cout());
defparam \ShiftRight0~121 .lut_mask = 16'hAACC;
defparam \ShiftRight0~121 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~122 (
	.dataa(csr_io_alu_op1_01),
	.datab(\_T_8~0_combout ),
	.datac(csr_io_alu_op2_01),
	.datad(csr_io_alu_op1_1),
	.cin(gnd),
	.combout(\ShiftRight0~122_combout ),
	.cout());
defparam \ShiftRight0~122 .lut_mask = 16'hF838;
defparam \ShiftRight0~122 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~123 (
	.dataa(alu_io_op1_31),
	.datab(alu_io_op1_30),
	.datac(\_T_8~0_combout ),
	.datad(\ShiftRight0~122_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~123_combout ),
	.cout());
defparam \ShiftRight0~123 .lut_mask = 16'hFC0A;
defparam \ShiftRight0~123 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~124 (
	.dataa(csr_io_alu_op2_11),
	.datab(alu_io_op2_210),
	.datac(\ShiftRight0~121_combout ),
	.datad(\ShiftRight0~123_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~124_combout ),
	.cout());
defparam \ShiftRight0~124 .lut_mask = 16'h5140;
defparam \ShiftRight0~124 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~125 (
	.dataa(\ShiftRight0~116_combout ),
	.datab(\ShiftRight0~120_combout ),
	.datac(\ShiftRight0~124_combout ),
	.datad(alu_io_op2_32),
	.cin(gnd),
	.combout(\ShiftRight0~125_combout ),
	.cout());
defparam \ShiftRight0~125 .lut_mask = 16'hAAFC;
defparam \ShiftRight0~125 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~127 (
	.dataa(csr_io_alu_op2_01),
	.datab(csr_io_alu_op2_11),
	.datac(alu_io_op2_32),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~127_combout ),
	.cout());
defparam \ShiftRight0~127 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~127 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[31]~47 (
	.dataa(csr_io_alu_op2_01),
	.datab(csr_io_alu_op1_02),
	.datac(ShiftRight02),
	.datad(ex_ctrl_alu_func_0),
	.cin(gnd),
	.combout(\op2_inv[31]~47_combout ),
	.cout());
defparam \op2_inv[31]~47 .lut_mask = 16'hF066;
defparam \op2_inv[31]~47 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[31]~43 (
	.dataa(ShiftRight03),
	.datab(_T_3_0),
	.datac(gnd),
	.datad(ex_ctrl_alu_func_0),
	.cin(gnd),
	.combout(\op2_inv[31]~43_combout ),
	.cout());
defparam \op2_inv[31]~43 .lut_mask = 16'hAACC;
defparam \op2_inv[31]~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[0]~0 (
	.dataa(ex_ctrl_alu_func_1),
	.datab(\op2_inv[31]~47_combout ),
	.datac(ex_ctrl_alu_func_2),
	.datad(\op2_inv[31]~43_combout ),
	.cin(gnd),
	.combout(\io_out[0]~0_combout ),
	.cout());
defparam \io_out[0]~0 .lut_mask = 16'hE5E0;
defparam \io_out[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \op2_inv[31]~44 (
	.dataa(csr_io_alu_op2_01),
	.datab(csr_io_alu_op1_02),
	.datac(gnd),
	.datad(ex_ctrl_alu_func_0),
	.cin(gnd),
	.combout(\op2_inv[31]~44_combout ),
	.cout());
defparam \op2_inv[31]~44 .lut_mask = 16'h88EE;
defparam \op2_inv[31]~44 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~129 (
	.dataa(alu_io_op2_32),
	.datab(alu_io_op2_210),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~129_combout ),
	.cout());
defparam \ShiftRight0~129 .lut_mask = 16'hEEEE;
defparam \ShiftRight0~129 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~131 (
	.dataa(\_T_60~combout ),
	.datab(csr_io_alu_op1_0),
	.datac(\ShiftRight0~34_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~131_combout ),
	.cout());
defparam \ShiftRight0~131 .lut_mask = 16'hAAC0;
defparam \ShiftRight0~131 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~132 (
	.dataa(\ShiftRight0~106_combout ),
	.datab(\ShiftRight0~103_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~132_combout ),
	.cout());
defparam \ShiftRight0~132 .lut_mask = 16'hAACC;
defparam \ShiftRight0~132 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~133 (
	.dataa(\ShiftRight0~131_combout ),
	.datab(csr_io_alu_op1_0),
	.datac(\ShiftRight0~132_combout ),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~133_combout ),
	.cout());
defparam \ShiftRight0~133 .lut_mask = 16'hAAC0;
defparam \ShiftRight0~133 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~134 (
	.dataa(csr_io_alu_op1_0),
	.datab(csr_io_alu_op2_11),
	.datac(csr_io_alu_op2_1),
	.datad(alu_io_op2_2),
	.cin(gnd),
	.combout(\ShiftRight0~134_combout ),
	.cout());
defparam \ShiftRight0~134 .lut_mask = 16'h0888;
defparam \ShiftRight0~134 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~135 (
	.dataa(csr_io_alu_op1_0),
	.datab(csr_io_alu_op2_1),
	.datac(alu_io_op2_2),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~135_combout ),
	.cout());
defparam \ShiftRight0~135 .lut_mask = 16'h002A;
defparam \ShiftRight0~135 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~136 (
	.dataa(\ShiftRight0~95_combout ),
	.datab(\ShiftRight0~100_combout ),
	.datac(\ShiftRight0~134_combout ),
	.datad(\ShiftRight0~135_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~136_combout ),
	.cout());
defparam \ShiftRight0~136 .lut_mask = 16'hEAC0;
defparam \ShiftRight0~136 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~137 (
	.dataa(csr_io_alu_op1_0),
	.datab(csr_io_alu_op2_11),
	.datac(alu_io_op2_210),
	.datad(\ShiftRight0~104_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~137_combout ),
	.cout());
defparam \ShiftRight0~137 .lut_mask = 16'h8000;
defparam \ShiftRight0~137 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~138 (
	.dataa(csr_io_alu_op1_0),
	.datab(csr_io_alu_op2_1),
	.datac(alu_io_op2_2),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~138_combout ),
	.cout());
defparam \ShiftRight0~138 .lut_mask = 16'h0080;
defparam \ShiftRight0~138 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~139 (
	.dataa(\ShiftRight0~136_combout ),
	.datab(\ShiftRight0~137_combout ),
	.datac(\ShiftRight0~99_combout ),
	.datad(\ShiftRight0~138_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~139_combout ),
	.cout());
defparam \ShiftRight0~139 .lut_mask = 16'hFEEE;
defparam \ShiftRight0~139 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~140 (
	.dataa(alu_io_op2_41),
	.datab(\ShiftRight0~133_combout ),
	.datac(\ShiftRight0~139_combout ),
	.datad(alu_io_op2_32),
	.cin(gnd),
	.combout(\ShiftRight0~140_combout ),
	.cout());
defparam \ShiftRight0~140 .lut_mask = 16'h88A0;
defparam \ShiftRight0~140 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~141 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~110_combout ),
	.datac(\ShiftRight0~117_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~141_combout ),
	.cout());
defparam \ShiftRight0~141 .lut_mask = 16'h88A0;
defparam \ShiftRight0~141 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~142 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~47_combout ),
	.datac(\ShiftRight0~42_combout ),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~142_combout ),
	.cout());
defparam \ShiftRight0~142 .lut_mask = 16'h88A0;
defparam \ShiftRight0~142 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~143 (
	.dataa(alu_io_op2_32),
	.datab(csr_io_alu_op2_11),
	.datac(gnd),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~143_combout ),
	.cout());
defparam \ShiftRight0~143 .lut_mask = 16'hAAEE;
defparam \ShiftRight0~143 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~144 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~118_combout ),
	.datac(csr_io_alu_op2_01),
	.datad(\ShiftRight0~43_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~144_combout ),
	.cout());
defparam \ShiftRight0~144 .lut_mask = 16'hA888;
defparam \ShiftRight0~144 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~145 (
	.dataa(\ShiftRight0~129_combout ),
	.datab(\ShiftRight0~142_combout ),
	.datac(\ShiftRight0~143_combout ),
	.datad(\ShiftRight0~144_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~145_combout ),
	.cout());
defparam \ShiftRight0~145 .lut_mask = 16'hE5E0;
defparam \ShiftRight0~145 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~146 (
	.dataa(\ShiftRight0~109_combout ),
	.datab(\ShiftRight0~114_combout ),
	.datac(\ShiftRight0~134_combout ),
	.datad(\ShiftRight0~135_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~146_combout ),
	.cout());
defparam \ShiftRight0~146 .lut_mask = 16'hEAC0;
defparam \ShiftRight0~146 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~147 (
	.dataa(csr_io_alu_op1_0),
	.datab(csr_io_alu_op2_11),
	.datac(alu_io_op2_210),
	.datad(\ShiftRight0~97_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~147_combout ),
	.cout());
defparam \ShiftRight0~147 .lut_mask = 16'h8000;
defparam \ShiftRight0~147 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~148 (
	.dataa(\ShiftRight0~146_combout ),
	.datab(\ShiftRight0~147_combout ),
	.datac(\ShiftRight0~113_combout ),
	.datad(\ShiftRight0~138_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~148_combout ),
	.cout());
defparam \ShiftRight0~148 .lut_mask = 16'hFEEE;
defparam \ShiftRight0~148 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~149 (
	.dataa(\ShiftRight0~141_combout ),
	.datab(\ShiftRight0~129_combout ),
	.datac(\ShiftRight0~145_combout ),
	.datad(\ShiftRight0~148_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~149_combout ),
	.cout());
defparam \ShiftRight0~149 .lut_mask = 16'hF838;
defparam \ShiftRight0~149 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~151 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~34_combout ),
	.datac(\ShiftRight0~106_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~151_combout ),
	.cout());
defparam \ShiftRight0~151 .lut_mask = 16'h88A0;
defparam \ShiftRight0~151 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~153 (
	.dataa(\ShiftRight0~69_combout ),
	.datab(\ShiftRight0~73_combout ),
	.datac(\ShiftRight0~135_combout ),
	.datad(\ShiftRight0~134_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~153_combout ),
	.cout());
defparam \ShiftRight0~153 .lut_mask = 16'hEAC0;
defparam \ShiftRight0~153 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~154 (
	.dataa(\_T_60~combout ),
	.datab(\_T_62[31]~0_combout ),
	.datac(csr_io_alu_op2_01),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~154_combout ),
	.cout());
defparam \ShiftRight0~154 .lut_mask = 16'hAAAC;
defparam \ShiftRight0~154 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~155 (
	.dataa(\ShiftRight0~153_combout ),
	.datab(alu_io_op2_210),
	.datac(\ShiftRight0~154_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~155_combout ),
	.cout());
defparam \ShiftRight0~155 .lut_mask = 16'hEAEA;
defparam \ShiftRight0~155 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~156 (
	.dataa(\ShiftRight0~91_combout ),
	.datab(\ShiftRight0~81_combout ),
	.datac(csr_io_alu_op2_11),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~156_combout ),
	.cout());
defparam \ShiftRight0~156 .lut_mask = 16'h00AC;
defparam \ShiftRight0~156 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~157 (
	.dataa(alu_io_op2_210),
	.datab(\ShiftRight0~76_combout ),
	.datac(\ShiftRight0~88_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~157_combout ),
	.cout());
defparam \ShiftRight0~157 .lut_mask = 16'h88A0;
defparam \ShiftRight0~157 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~244 (
	.dataa(ex_ctrl_alu_op1_0),
	.datab(ex_ctrl_alu_op1_1),
	.datac(\ShiftRight0~156_combout ),
	.datad(\ShiftRight0~157_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~244_combout ),
	.cout());
defparam \ShiftRight0~244 .lut_mask = 16'h6660;
defparam \ShiftRight0~244 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~158 (
	.dataa(alu_io_op2_41),
	.datab(\ShiftRight0~155_combout ),
	.datac(\ShiftRight0~244_combout ),
	.datad(alu_io_op2_32),
	.cin(gnd),
	.combout(\ShiftRight0~158_combout ),
	.cout());
defparam \ShiftRight0~158 .lut_mask = 16'h88A0;
defparam \ShiftRight0~158 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~159 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~46_combout ),
	.datac(\ShiftRight0~47_combout ),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~159_combout ),
	.cout());
defparam \ShiftRight0~159 .lut_mask = 16'h88A0;
defparam \ShiftRight0~159 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~160 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~58_combout ),
	.datac(\ShiftRight0~41_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~160_combout ),
	.cout());
defparam \ShiftRight0~160 .lut_mask = 16'h88A0;
defparam \ShiftRight0~160 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~161 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~42_combout ),
	.datac(\ShiftRight0~43_combout ),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~161_combout ),
	.cout());
defparam \ShiftRight0~161 .lut_mask = 16'h88A0;
defparam \ShiftRight0~161 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~162 (
	.dataa(\ShiftRight0~143_combout ),
	.datab(\ShiftRight0~160_combout ),
	.datac(\ShiftRight0~129_combout ),
	.datad(\ShiftRight0~161_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~162_combout ),
	.cout());
defparam \ShiftRight0~162 .lut_mask = 16'hE5E0;
defparam \ShiftRight0~162 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~163 (
	.dataa(\ShiftRight0~84_combout ),
	.datab(\ShiftRight0~60_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~163_combout ),
	.cout());
defparam \ShiftRight0~163 .lut_mask = 16'hAACC;
defparam \ShiftRight0~163 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~164 (
	.dataa(\ShiftRight0~63_combout ),
	.datab(\ShiftRight0~55_combout ),
	.datac(gnd),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~164_combout ),
	.cout());
defparam \ShiftRight0~164 .lut_mask = 16'hAACC;
defparam \ShiftRight0~164 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~165 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~163_combout ),
	.datac(\ShiftRight0~164_combout ),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~165_combout ),
	.cout());
defparam \ShiftRight0~165 .lut_mask = 16'h88A0;
defparam \ShiftRight0~165 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~166 (
	.dataa(\ShiftRight0~159_combout ),
	.datab(\ShiftRight0~143_combout ),
	.datac(\ShiftRight0~162_combout ),
	.datad(\ShiftRight0~165_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~166_combout ),
	.cout());
defparam \ShiftRight0~166 .lut_mask = 16'hF838;
defparam \ShiftRight0~166 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~168 (
	.dataa(gnd),
	.datab(csr_io_alu_op2_1),
	.datac(alu_io_op2_2),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~168_combout ),
	.cout());
defparam \ShiftRight0~168 .lut_mask = 16'h003F;
defparam \ShiftRight0~168 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~169 (
	.dataa(\_T_60~combout ),
	.datab(\_T_62[31]~0_combout ),
	.datac(\ShiftRight0~168_combout ),
	.datad(csr_io_alu_op2_01),
	.cin(gnd),
	.combout(\ShiftRight0~169_combout ),
	.cout());
defparam \ShiftRight0~169 .lut_mask = 16'hAACA;
defparam \ShiftRight0~169 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~170 (
	.dataa(csr_io_alu_op2_11),
	.datab(alu_io_op2_210),
	.datac(\ShiftRight0~69_combout ),
	.datad(\ShiftRight0~73_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~170_combout ),
	.cout());
defparam \ShiftRight0~170 .lut_mask = 16'hE6A2;
defparam \ShiftRight0~170 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~171 (
	.dataa(\ShiftRight0~76_combout ),
	.datab(\ShiftRight0~88_combout ),
	.datac(alu_io_op2_210),
	.datad(\ShiftRight0~170_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~171_combout ),
	.cout());
defparam \ShiftRight0~171 .lut_mask = 16'hFA0C;
defparam \ShiftRight0~171 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~172 (
	.dataa(\ShiftRight0~169_combout ),
	.datab(csr_io_alu_op1_0),
	.datac(\ShiftRight0~171_combout ),
	.datad(alu_io_op2_32),
	.cin(gnd),
	.combout(\ShiftRight0~172_combout ),
	.cout());
defparam \ShiftRight0~172 .lut_mask = 16'hAAC0;
defparam \ShiftRight0~172 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~245 (
	.dataa(ex_ctrl_alu_op1_0),
	.datab(ex_ctrl_alu_op1_1),
	.datac(\ShiftRight0~105_combout ),
	.datad(\ShiftRight0~107_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~245_combout ),
	.cout());
defparam \ShiftRight0~245 .lut_mask = 16'h6660;
defparam \ShiftRight0~245 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~246 (
	.dataa(ex_ctrl_alu_op1_0),
	.datab(ex_ctrl_alu_op1_1),
	.datac(\ShiftRight0~98_combout ),
	.datad(\ShiftRight0~101_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~246_combout ),
	.cout());
defparam \ShiftRight0~246 .lut_mask = 16'h6660;
defparam \ShiftRight0~246 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~247 (
	.dataa(ex_ctrl_alu_op1_0),
	.datab(ex_ctrl_alu_op1_1),
	.datac(\ShiftRight0~111_combout ),
	.datad(\ShiftRight0~115_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~247_combout ),
	.cout());
defparam \ShiftRight0~247 .lut_mask = 16'h6660;
defparam \ShiftRight0~247 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~174 (
	.dataa(alu_io_op2_41),
	.datab(\ShiftRight0~246_combout ),
	.datac(alu_io_op2_32),
	.datad(\ShiftRight0~247_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~174_combout ),
	.cout());
defparam \ShiftRight0~174 .lut_mask = 16'hE5E0;
defparam \ShiftRight0~174 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~176 (
	.dataa(\_T_60~combout ),
	.datab(csr_io_alu_op1_0),
	.datac(\ShiftRight0~34_combout ),
	.datad(\ShiftRight0~242_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~176_combout ),
	.cout());
defparam \ShiftRight0~176 .lut_mask = 16'hAAC0;
defparam \ShiftRight0~176 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~177 (
	.dataa(csr_io_alu_op2_11),
	.datab(alu_io_op2_210),
	.datac(\ShiftRight0~106_combout ),
	.datad(\ShiftRight0~103_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~177_combout ),
	.cout());
defparam \ShiftRight0~177 .lut_mask = 16'hE6A2;
defparam \ShiftRight0~177 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~178 (
	.dataa(\ShiftRight0~104_combout ),
	.datab(\ShiftRight0~99_combout ),
	.datac(alu_io_op2_210),
	.datad(\ShiftRight0~177_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~178_combout ),
	.cout());
defparam \ShiftRight0~178 .lut_mask = 16'hFA0C;
defparam \ShiftRight0~178 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~179 (
	.dataa(\ShiftRight0~176_combout ),
	.datab(csr_io_alu_op1_0),
	.datac(\ShiftRight0~178_combout ),
	.datad(alu_io_op2_32),
	.cin(gnd),
	.combout(\ShiftRight0~179_combout ),
	.cout());
defparam \ShiftRight0~179 .lut_mask = 16'hAAC0;
defparam \ShiftRight0~179 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~181 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~59_combout ),
	.datac(alu_io_op2_210),
	.datad(\ShiftRight0~64_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~181_combout ),
	.cout());
defparam \ShiftRight0~181 .lut_mask = 16'hA888;
defparam \ShiftRight0~181 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~182 (
	.dataa(alu_io_op2_32),
	.datab(\ShiftRight0~78_combout ),
	.datac(alu_io_op2_41),
	.datad(\ShiftRight0~181_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~182_combout ),
	.cout());
defparam \ShiftRight0~182 .lut_mask = 16'hE5E0;
defparam \ShiftRight0~182 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~184 (
	.dataa(alu_io_op2_32),
	.datab(\_T_60~combout ),
	.datac(\ShiftRight0~70_combout ),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~184_combout ),
	.cout());
defparam \ShiftRight0~184 .lut_mask = 16'h88A0;
defparam \ShiftRight0~184 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~185 (
	.dataa(csr_io_alu_op2_11),
	.datab(alu_io_op2_210),
	.datac(\ShiftRight0~73_combout ),
	.datad(\ShiftRight0~76_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~185_combout ),
	.cout());
defparam \ShiftRight0~185 .lut_mask = 16'hE6A2;
defparam \ShiftRight0~185 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~186 (
	.dataa(\ShiftRight0~88_combout ),
	.datab(\ShiftRight0~91_combout ),
	.datac(alu_io_op2_210),
	.datad(\ShiftRight0~185_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~186_combout ),
	.cout());
defparam \ShiftRight0~186 .lut_mask = 16'hFA0C;
defparam \ShiftRight0~186 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~187 (
	.dataa(\ShiftRight0~184_combout ),
	.datab(csr_io_alu_op1_0),
	.datac(\ShiftRight0~186_combout ),
	.datad(alu_io_op2_32),
	.cin(gnd),
	.combout(\ShiftRight0~187_combout ),
	.cout());
defparam \ShiftRight0~187 .lut_mask = 16'hAAEA;
defparam \ShiftRight0~187 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~189 (
	.dataa(alu_io_op2_41),
	.datab(\ShiftRight0~139_combout ),
	.datac(alu_io_op2_32),
	.datad(\ShiftRight0~148_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~189_combout ),
	.cout());
defparam \ShiftRight0~189 .lut_mask = 16'hE5E0;
defparam \ShiftRight0~189 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~191 (
	.dataa(alu_io_op2_32),
	.datab(\_T_60~combout ),
	.datac(\ShiftRight0~151_combout ),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~191_combout ),
	.cout());
defparam \ShiftRight0~191 .lut_mask = 16'h88A0;
defparam \ShiftRight0~191 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~192 (
	.dataa(csr_io_alu_op2_11),
	.datab(alu_io_op2_210),
	.datac(\ShiftRight0~103_combout ),
	.datad(\ShiftRight0~104_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~192_combout ),
	.cout());
defparam \ShiftRight0~192 .lut_mask = 16'hE6A2;
defparam \ShiftRight0~192 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~193 (
	.dataa(\ShiftRight0~99_combout ),
	.datab(\ShiftRight0~100_combout ),
	.datac(alu_io_op2_210),
	.datad(\ShiftRight0~192_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~193_combout ),
	.cout());
defparam \ShiftRight0~193 .lut_mask = 16'hFA0C;
defparam \ShiftRight0~193 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~194 (
	.dataa(\ShiftRight0~191_combout ),
	.datab(csr_io_alu_op1_0),
	.datac(\ShiftRight0~193_combout ),
	.datad(alu_io_op2_32),
	.cin(gnd),
	.combout(\ShiftRight0~194_combout ),
	.cout());
defparam \ShiftRight0~194 .lut_mask = 16'hAAEA;
defparam \ShiftRight0~194 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~196 (
	.dataa(alu_io_op2_32),
	.datab(\ShiftRight0~155_combout ),
	.datac(alu_io_op2_41),
	.datad(\ShiftRight0~165_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~196_combout ),
	.cout());
defparam \ShiftRight0~196 .lut_mask = 16'hE5E0;
defparam \ShiftRight0~196 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~248 (
	.dataa(alu_io_op2_32),
	.datab(alu_io_op2_41),
	.datac(\ShiftRight0~244_combout ),
	.datad(\_T_60~combout ),
	.cin(gnd),
	.combout(\ShiftRight0~248_combout ),
	.cout());
defparam \ShiftRight0~248 .lut_mask = 16'hDC10;
defparam \ShiftRight0~248 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~199 (
	.dataa(alu_io_op2_41),
	.datab(\_T_60~combout ),
	.datac(\ShiftRight0~151_combout ),
	.datad(\ShiftRight0~129_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~199_combout ),
	.cout());
defparam \ShiftRight0~199 .lut_mask = 16'h88A0;
defparam \ShiftRight0~199 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~200 (
	.dataa(\ShiftRight0~113_combout ),
	.datab(\ShiftRight0~114_combout ),
	.datac(csr_io_alu_op2_11),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~200_combout ),
	.cout());
defparam \ShiftRight0~200 .lut_mask = 16'h00AC;
defparam \ShiftRight0~200 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~201 (
	.dataa(alu_io_op2_210),
	.datab(\ShiftRight0~95_combout ),
	.datac(\ShiftRight0~97_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~201_combout ),
	.cout());
defparam \ShiftRight0~201 .lut_mask = 16'h88A0;
defparam \ShiftRight0~201 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~202 (
	.dataa(\ShiftRight0~200_combout ),
	.datab(\ShiftRight0~201_combout ),
	.datac(\ShiftRight0~193_combout ),
	.datad(alu_io_op2_32),
	.cin(gnd),
	.combout(\ShiftRight0~202_combout ),
	.cout());
defparam \ShiftRight0~202 .lut_mask = 16'hF0EE;
defparam \ShiftRight0~202 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~205 (
	.dataa(alu_io_op2_41),
	.datab(\_T_60~combout ),
	.datac(\ShiftRight0~70_combout ),
	.datad(\ShiftRight0~129_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~205_combout ),
	.cout());
defparam \ShiftRight0~205 .lut_mask = 16'h88A0;
defparam \ShiftRight0~205 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~206 (
	.dataa(alu_io_op2_210),
	.datab(\ShiftRight0~81_combout ),
	.datac(\ShiftRight0~84_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~206_combout ),
	.cout());
defparam \ShiftRight0~206 .lut_mask = 16'h88A0;
defparam \ShiftRight0~206 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~207 (
	.dataa(\ShiftRight0~206_combout ),
	.datab(\ShiftRight0~64_combout ),
	.datac(gnd),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~207_combout ),
	.cout());
defparam \ShiftRight0~207 .lut_mask = 16'hAAEE;
defparam \ShiftRight0~207 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~208 (
	.dataa(\ShiftRight0~241_combout ),
	.datab(\ShiftRight0~186_combout ),
	.datac(\ShiftRight0~207_combout ),
	.datad(alu_io_op2_32),
	.cin(gnd),
	.combout(\ShiftRight0~208_combout ),
	.cout());
defparam \ShiftRight0~208 .lut_mask = 16'h88A0;
defparam \ShiftRight0~208 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~211 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~34_combout ),
	.datac(\ShiftRight0~242_combout ),
	.datad(\_T_60~combout ),
	.cin(gnd),
	.combout(\ShiftRight0~211_combout ),
	.cout());
defparam \ShiftRight0~211 .lut_mask = 16'hF808;
defparam \ShiftRight0~211 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~212 (
	.dataa(alu_io_op2_32),
	.datab(alu_io_op2_41),
	.datac(\_T_60~combout ),
	.datad(\ShiftRight0~211_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~212_combout ),
	.cout());
defparam \ShiftRight0~212 .lut_mask = 16'hC480;
defparam \ShiftRight0~212 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~213 (
	.dataa(\ShiftRight0~97_combout ),
	.datab(\ShiftRight0~113_combout ),
	.datac(csr_io_alu_op2_11),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~213_combout ),
	.cout());
defparam \ShiftRight0~213 .lut_mask = 16'h00AC;
defparam \ShiftRight0~213 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~214 (
	.dataa(alu_io_op2_210),
	.datab(\ShiftRight0~100_combout ),
	.datac(\ShiftRight0~95_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~214_combout ),
	.cout());
defparam \ShiftRight0~214 .lut_mask = 16'h88A0;
defparam \ShiftRight0~214 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~215 (
	.dataa(\ShiftRight0~213_combout ),
	.datab(\ShiftRight0~214_combout ),
	.datac(\ShiftRight0~178_combout ),
	.datad(alu_io_op2_32),
	.cin(gnd),
	.combout(\ShiftRight0~215_combout ),
	.cout());
defparam \ShiftRight0~215 .lut_mask = 16'hF0EE;
defparam \ShiftRight0~215 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~218 (
	.dataa(alu_io_op2_41),
	.datab(\_T_60~combout ),
	.datac(\_T_62[31]~0_combout ),
	.datad(\ShiftRight0~127_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~218_combout ),
	.cout());
defparam \ShiftRight0~218 .lut_mask = 16'h88A0;
defparam \ShiftRight0~218 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~219 (
	.dataa(alu_io_op2_210),
	.datab(\ShiftRight0~91_combout ),
	.datac(\ShiftRight0~81_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~219_combout ),
	.cout());
defparam \ShiftRight0~219 .lut_mask = 16'h88A0;
defparam \ShiftRight0~219 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~220 (
	.dataa(\ShiftRight0~219_combout ),
	.datab(\ShiftRight0~163_combout ),
	.datac(gnd),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~220_combout ),
	.cout());
defparam \ShiftRight0~220 .lut_mask = 16'hAAEE;
defparam \ShiftRight0~220 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~221 (
	.dataa(\ShiftRight0~241_combout ),
	.datab(\ShiftRight0~171_combout ),
	.datac(\ShiftRight0~220_combout ),
	.datad(alu_io_op2_32),
	.cin(gnd),
	.combout(\ShiftRight0~221_combout ),
	.cout());
defparam \ShiftRight0~221 .lut_mask = 16'h88A0;
defparam \ShiftRight0~221 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~223 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~109_combout ),
	.datac(\ShiftRight0~110_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~223_combout ),
	.cout());
defparam \ShiftRight0~223 .lut_mask = 16'h88A0;
defparam \ShiftRight0~223 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~224 (
	.dataa(alu_io_op2_4),
	.datab(io_sw_r_ex_imm_4),
	.datac(ex_ctrl_alu_op210),
	.datad(\ShiftRight0~37_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~224_combout ),
	.cout());
defparam \ShiftRight0~224 .lut_mask = 16'h00AE;
defparam \ShiftRight0~224 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~225 (
	.dataa(csr_io_alu_op2_1),
	.datab(\ShiftRight0~224_combout ),
	.datac(alu_io_op2_2),
	.datad(\ShiftRight0~37_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~225_combout ),
	.cout());
defparam \ShiftRight0~225 .lut_mask = 16'hA888;
defparam \ShiftRight0~225 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~252 (
	.dataa(ex_ctrl_alu_op1_0),
	.datab(ex_ctrl_alu_op1_1),
	.datac(\ShiftRight0~200_combout ),
	.datad(\ShiftRight0~201_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~252_combout ),
	.cout());
defparam \ShiftRight0~252 .lut_mask = 16'h6660;
defparam \ShiftRight0~252 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~226 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~117_combout ),
	.datac(\ShiftRight0~121_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~226_combout ),
	.cout());
defparam \ShiftRight0~226 .lut_mask = 16'h88A0;
defparam \ShiftRight0~226 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~227 (
	.dataa(\ShiftRight0~225_combout ),
	.datab(\ShiftRight0~252_combout ),
	.datac(\ShiftRight0~37_combout ),
	.datad(\ShiftRight0~226_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~227_combout ),
	.cout());
defparam \ShiftRight0~227 .lut_mask = 16'h5E0E;
defparam \ShiftRight0~227 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~229 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~206_combout ),
	.datac(\ShiftRight0~64_combout ),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~229_combout ),
	.cout());
defparam \ShiftRight0~229 .lut_mask = 16'h88A8;
defparam \ShiftRight0~229 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~230 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~55_combout ),
	.datac(\ShiftRight0~58_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~230_combout ),
	.cout());
defparam \ShiftRight0~230 .lut_mask = 16'h88A0;
defparam \ShiftRight0~230 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~231 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~41_combout ),
	.datac(\ShiftRight0~48_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~231_combout ),
	.cout());
defparam \ShiftRight0~231 .lut_mask = 16'h88A0;
defparam \ShiftRight0~231 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~232 (
	.dataa(\ShiftRight0~37_combout ),
	.datab(\ShiftRight0~230_combout ),
	.datac(\ShiftRight0~225_combout ),
	.datad(\ShiftRight0~231_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~232_combout ),
	.cout());
defparam \ShiftRight0~232 .lut_mask = 16'hDAD0;
defparam \ShiftRight0~232 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~234 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~114_combout ),
	.datac(\ShiftRight0~109_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~234_combout ),
	.cout());
defparam \ShiftRight0~234 .lut_mask = 16'h88A0;
defparam \ShiftRight0~234 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~255 (
	.dataa(ex_ctrl_alu_op1_0),
	.datab(ex_ctrl_alu_op1_1),
	.datac(\ShiftRight0~213_combout ),
	.datad(\ShiftRight0~214_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~255_combout ),
	.cout());
defparam \ShiftRight0~255 .lut_mask = 16'h6660;
defparam \ShiftRight0~255 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~235 (
	.dataa(\ShiftRight0~225_combout ),
	.datab(\ShiftRight0~255_combout ),
	.datac(\ShiftRight0~37_combout ),
	.datad(\ShiftRight0~141_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~235_combout ),
	.cout());
defparam \ShiftRight0~235 .lut_mask = 16'h5E0E;
defparam \ShiftRight0~235 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~237 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~219_combout ),
	.datac(\ShiftRight0~163_combout ),
	.datad(alu_io_op2_210),
	.cin(gnd),
	.combout(\ShiftRight0~237_combout ),
	.cout());
defparam \ShiftRight0~237 .lut_mask = 16'h88A8;
defparam \ShiftRight0~237 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~238 (
	.dataa(csr_io_alu_op1_0),
	.datab(\ShiftRight0~63_combout ),
	.datac(\ShiftRight0~55_combout ),
	.datad(csr_io_alu_op2_11),
	.cin(gnd),
	.combout(\ShiftRight0~238_combout ),
	.cout());
defparam \ShiftRight0~238 .lut_mask = 16'h88A0;
defparam \ShiftRight0~238 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~239 (
	.dataa(\ShiftRight0~37_combout ),
	.datab(\ShiftRight0~238_combout ),
	.datac(\ShiftRight0~225_combout ),
	.datad(\ShiftRight0~160_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~239_combout ),
	.cout());
defparam \ShiftRight0~239 .lut_mask = 16'hDAD0;
defparam \ShiftRight0~239 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~204 (
	.dataa(\_T_60~combout ),
	.datab(alu_io_op2_32),
	.datac(\ShiftRight0~133_combout ),
	.datad(alu_io_op2_41),
	.cin(gnd),
	.combout(\ShiftRight0~204_combout ),
	.cout());
defparam \ShiftRight0~204 .lut_mask = 16'hAAC0;
defparam \ShiftRight0~204 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \ShiftRight0~210 (
	.dataa(\_T_60~combout ),
	.datab(alu_io_op2_32),
	.datac(\ShiftRight0~78_combout ),
	.datad(alu_io_op2_41),
	.cin(gnd),
	.combout(\ShiftRight0~210_combout ),
	.cout());
defparam \ShiftRight0~210 .lut_mask = 16'hAAC0;
defparam \ShiftRight0~210 .sum_lutc_input = "datac";

endmodule

module kyogenrv_fpga_CSR (
	ex_j_check,
	ex_ctrl_mem_wr01,
	_T_3549,
	mepc_2,
	mepc_3,
	mepc_4,
	mepc_5,
	mepc_6,
	mepc_7,
	mepc_8,
	mepc_9,
	mepc_10,
	mepc_11,
	mepc_12,
	mepc_13,
	mepc_14,
	mepc_15,
	mepc_16,
	mepc_17,
	mepc_18,
	mepc_19,
	mepc_20,
	mepc_21,
	mepc_22,
	mepc_23,
	mepc_24,
	mepc_25,
	mepc_26,
	mepc_27,
	mepc_28,
	mepc_29,
	mepc_30,
	mepc_31,
	ex_b_check,
	inst_kill,
	ex_npc_0,
	ex_npc_1,
	Equal56,
	ex_pc_4,
	ex_pc_5,
	ex_pc_6,
	ex_pc_7,
	ex_pc_2,
	ex_pc_3,
	ex_pc_8,
	ex_pc_9,
	ex_pc_10,
	ex_pc_11,
	ex_pc_12,
	ex_pc_13,
	ex_pc_14,
	ex_pc_15,
	ex_pc_16,
	ex_pc_17,
	ex_pc_18,
	ex_pc_19,
	ex_pc_20,
	ex_pc_21,
	ex_pc_22,
	ex_pc_23,
	ex_pc_24,
	ex_pc_25,
	ex_pc_26,
	ex_pc_27,
	ex_pc_28,
	ex_pc_29,
	ex_pc_30,
	ex_pc_31,
	Equal561,
	ex_ctrl_legal,
	Equal59,
	ex_csr_addr_0,
	ex_csr_addr_1,
	ex_csr_addr_2,
	ex_csr_addr_3,
	ex_csr_addr_4,
	Equal62,
	ex_inst_8,
	ex_ctrl_imm_type001,
	csr_io_alu_op2_1,
	ex_inst_7,
	csr_io_alu_op2_0,
	ex_ctrl_mask_type_0,
	ex_ctrl_mask_type_2,
	ex_ctrl_mask_type_1,
	io_expt1,
	waitrequest_reset_override,
	wait_latency_counter_0,
	mem_ctrl_mem_wr10,
	wait_latency_counter_1,
	read_latency_shift_reg_0,
	ex_inst_9,
	ex_inst_10,
	ex_inst_11,
	_T_3557,
	mcause_0,
	ex_csr_cmd_2,
	ex_csr_cmd_0,
	ex_csr_cmd_1,
	ex_csr_addr_8,
	isEcall,
	altera_reset_synchronizer_int_chain_out,
	mepc_0,
	io_expt2,
	mtvec_0,
	ex_csr_addr_9,
	ex_csr_addr_11,
	ex_csr_addr_10,
	ex_inst_13,
	ex_inst_12,
	ex_inst_14,
	ex_csr_addr_5,
	ex_csr_addr_6,
	ex_csr_addr_7,
	mepc_1,
	mtvec_1,
	io_out_1,
	io_out_0,
	mtvec_2,
	mtvec_3,
	mtvec_4,
	mtvec_5,
	mtvec_6,
	mtvec_7,
	mtvec_8,
	mtvec_9,
	mtvec_10,
	mtvec_11,
	mtvec_12,
	mtvec_13,
	mtvec_14,
	mtvec_15,
	mtvec_16,
	mtvec_17,
	mtvec_18,
	mtvec_19,
	mtvec_20,
	mtvec_21,
	mtvec_22,
	mtvec_23,
	mtvec_24,
	mtvec_25,
	mtvec_26,
	mtvec_27,
	mtvec_28,
	mtvec_29,
	mtvec_30,
	mtvec_31,
	csr_io_in_0,
	io_out_28,
	io_out_29,
	io_out_291,
	io_out_30,
	io_out_31,
	io_out_8,
	io_out_9,
	io_out_10,
	io_out_11,
	io_out_12,
	io_out_13,
	io_out_14,
	io_out_15,
	io_out_16,
	io_out_17,
	io_out_18,
	io_out_19,
	io_out_4,
	io_out_2,
	io_out_3,
	io_out_5,
	io_out_6,
	io_out_7,
	io_out_20,
	io_out_21,
	io_out_211,
	io_out_22,
	io_out_23,
	io_out_24,
	io_out_25,
	io_out_251,
	io_out_26,
	io_out_27,
	io_out_271,
	csr_io_in_1,
	ex_inst_0,
	ex_inst_1,
	ex_inst_4,
	ex_inst_2,
	ex_inst_3,
	ex_inst_5,
	ex_inst_6,
	csr_io_in_2,
	csr_io_in_3,
	csr_io_in_4,
	csr_io_in_5,
	csr_io_in_6,
	csr_io_in_7,
	csr_io_in_8,
	csr_io_in_9,
	csr_io_in_10,
	csr_io_in_11,
	csr_io_in_12,
	csr_io_in_13,
	csr_io_in_14,
	csr_io_in_15,
	csr_io_in_16,
	csr_io_in_17,
	csr_io_in_18,
	csr_io_in_19,
	csr_io_in_20,
	csr_io_in_21,
	csr_io_in_22,
	csr_io_in_23,
	csr_io_in_24,
	csr_io_in_25,
	csr_io_in_26,
	csr_io_in_27,
	csr_io_in_28,
	csr_io_in_29,
	csr_io_in_30,
	csr_io_in_31,
	csr_io_alu_op1_1,
	csr_io_alu_op1_0,
	clock)/* synthesis synthesis_greybox=0 */;
input 	ex_j_check;
input 	ex_ctrl_mem_wr01;
input 	_T_3549;
output 	mepc_2;
output 	mepc_3;
output 	mepc_4;
output 	mepc_5;
output 	mepc_6;
output 	mepc_7;
output 	mepc_8;
output 	mepc_9;
output 	mepc_10;
output 	mepc_11;
output 	mepc_12;
output 	mepc_13;
output 	mepc_14;
output 	mepc_15;
output 	mepc_16;
output 	mepc_17;
output 	mepc_18;
output 	mepc_19;
output 	mepc_20;
output 	mepc_21;
output 	mepc_22;
output 	mepc_23;
output 	mepc_24;
output 	mepc_25;
output 	mepc_26;
output 	mepc_27;
output 	mepc_28;
output 	mepc_29;
output 	mepc_30;
output 	mepc_31;
input 	ex_b_check;
input 	inst_kill;
input 	ex_npc_0;
input 	ex_npc_1;
input 	Equal56;
input 	ex_pc_4;
input 	ex_pc_5;
input 	ex_pc_6;
input 	ex_pc_7;
input 	ex_pc_2;
input 	ex_pc_3;
input 	ex_pc_8;
input 	ex_pc_9;
input 	ex_pc_10;
input 	ex_pc_11;
input 	ex_pc_12;
input 	ex_pc_13;
input 	ex_pc_14;
input 	ex_pc_15;
input 	ex_pc_16;
input 	ex_pc_17;
input 	ex_pc_18;
input 	ex_pc_19;
input 	ex_pc_20;
input 	ex_pc_21;
input 	ex_pc_22;
input 	ex_pc_23;
input 	ex_pc_24;
input 	ex_pc_25;
input 	ex_pc_26;
input 	ex_pc_27;
input 	ex_pc_28;
input 	ex_pc_29;
input 	ex_pc_30;
input 	ex_pc_31;
input 	Equal561;
input 	ex_ctrl_legal;
input 	Equal59;
input 	ex_csr_addr_0;
input 	ex_csr_addr_1;
input 	ex_csr_addr_2;
input 	ex_csr_addr_3;
input 	ex_csr_addr_4;
input 	Equal62;
input 	ex_inst_8;
input 	ex_ctrl_imm_type001;
input 	csr_io_alu_op2_1;
input 	ex_inst_7;
input 	csr_io_alu_op2_0;
input 	ex_ctrl_mask_type_0;
input 	ex_ctrl_mask_type_2;
input 	ex_ctrl_mask_type_1;
output 	io_expt1;
input 	waitrequest_reset_override;
input 	wait_latency_counter_0;
input 	mem_ctrl_mem_wr10;
input 	wait_latency_counter_1;
input 	read_latency_shift_reg_0;
input 	ex_inst_9;
input 	ex_inst_10;
input 	ex_inst_11;
input 	_T_3557;
output 	mcause_0;
input 	ex_csr_cmd_2;
input 	ex_csr_cmd_0;
input 	ex_csr_cmd_1;
input 	ex_csr_addr_8;
output 	isEcall;
input 	altera_reset_synchronizer_int_chain_out;
output 	mepc_0;
output 	io_expt2;
output 	mtvec_0;
input 	ex_csr_addr_9;
input 	ex_csr_addr_11;
input 	ex_csr_addr_10;
input 	ex_inst_13;
input 	ex_inst_12;
input 	ex_inst_14;
input 	ex_csr_addr_5;
input 	ex_csr_addr_6;
input 	ex_csr_addr_7;
output 	mepc_1;
output 	mtvec_1;
output 	io_out_1;
output 	io_out_0;
output 	mtvec_2;
output 	mtvec_3;
output 	mtvec_4;
output 	mtvec_5;
output 	mtvec_6;
output 	mtvec_7;
output 	mtvec_8;
output 	mtvec_9;
output 	mtvec_10;
output 	mtvec_11;
output 	mtvec_12;
output 	mtvec_13;
output 	mtvec_14;
output 	mtvec_15;
output 	mtvec_16;
output 	mtvec_17;
output 	mtvec_18;
output 	mtvec_19;
output 	mtvec_20;
output 	mtvec_21;
output 	mtvec_22;
output 	mtvec_23;
output 	mtvec_24;
output 	mtvec_25;
output 	mtvec_26;
output 	mtvec_27;
output 	mtvec_28;
output 	mtvec_29;
output 	mtvec_30;
output 	mtvec_31;
input 	csr_io_in_0;
output 	io_out_28;
output 	io_out_29;
output 	io_out_291;
output 	io_out_30;
output 	io_out_31;
output 	io_out_8;
output 	io_out_9;
output 	io_out_10;
output 	io_out_11;
output 	io_out_12;
output 	io_out_13;
output 	io_out_14;
output 	io_out_15;
output 	io_out_16;
output 	io_out_17;
output 	io_out_18;
output 	io_out_19;
output 	io_out_4;
output 	io_out_2;
output 	io_out_3;
output 	io_out_5;
output 	io_out_6;
output 	io_out_7;
output 	io_out_20;
output 	io_out_21;
output 	io_out_211;
output 	io_out_22;
output 	io_out_23;
output 	io_out_24;
output 	io_out_25;
output 	io_out_251;
output 	io_out_26;
output 	io_out_27;
output 	io_out_271;
input 	csr_io_in_1;
input 	ex_inst_0;
input 	ex_inst_1;
input 	ex_inst_4;
input 	ex_inst_2;
input 	ex_inst_3;
input 	ex_inst_5;
input 	ex_inst_6;
input 	csr_io_in_2;
input 	csr_io_in_3;
input 	csr_io_in_4;
input 	csr_io_in_5;
input 	csr_io_in_6;
input 	csr_io_in_7;
input 	csr_io_in_8;
input 	csr_io_in_9;
input 	csr_io_in_10;
input 	csr_io_in_11;
input 	csr_io_in_12;
input 	csr_io_in_13;
input 	csr_io_in_14;
input 	csr_io_in_15;
input 	csr_io_in_16;
input 	csr_io_in_17;
input 	csr_io_in_18;
input 	csr_io_in_19;
input 	csr_io_in_20;
input 	csr_io_in_21;
input 	csr_io_in_22;
input 	csr_io_in_23;
input 	csr_io_in_24;
input 	csr_io_in_25;
input 	csr_io_in_26;
input 	csr_io_in_27;
input 	csr_io_in_28;
input 	csr_io_in_29;
input 	csr_io_in_30;
input 	csr_io_in_31;
input 	csr_io_alu_op1_1;
input 	csr_io_alu_op1_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \pre_mepc~3_combout ;
wire \pre_mepc[28]~1_combout ;
wire \pre_mepc[2]~q ;
wire \mepc[2]~0_combout ;
wire \_T_246[0]~0_combout ;
wire \_T_246[2]~5_combout ;
wire \_T_246[2]~6_combout ;
wire \Equal19~0_combout ;
wire \Equal25~2_combout ;
wire \Equal16~0_combout ;
wire \Equal4~0_combout ;
wire \Equal26~0_combout ;
wire \wen~combout ;
wire \mepc[0]~30_combout ;
wire \pre_mepc~4_combout ;
wire \pre_mepc[3]~q ;
wire \mepc[3]~1_combout ;
wire \_T_246[3]~7_combout ;
wire \_T_246[3]~8_combout ;
wire \pre_mepc~5_combout ;
wire \pre_mepc[4]~q ;
wire \mepc[4]~2_combout ;
wire \_T_244[4]~0_combout ;
wire \_T_244[4]~1_combout ;
wire \pre_mepc~6_combout ;
wire \pre_mepc[5]~q ;
wire \mepc[5]~3_combout ;
wire \_T_244[5]~2_combout ;
wire \_T_244[5]~3_combout ;
wire \pre_mepc~7_combout ;
wire \pre_mepc[6]~q ;
wire \mepc[6]~4_combout ;
wire \_T_244[6]~4_combout ;
wire \_T_244[6]~5_combout ;
wire \pre_mepc~8_combout ;
wire \pre_mepc[7]~q ;
wire \mepc[7]~5_combout ;
wire \_T_244[7]~6_combout ;
wire \_T_244[7]~7_combout ;
wire \pre_mepc~9_combout ;
wire \pre_mepc[8]~q ;
wire \mepc[8]~6_combout ;
wire \_T_244[8]~8_combout ;
wire \_T_244[8]~9_combout ;
wire \pre_mepc~10_combout ;
wire \pre_mepc[9]~q ;
wire \mepc[9]~7_combout ;
wire \_T_244[9]~10_combout ;
wire \_T_244[9]~11_combout ;
wire \pre_mepc~11_combout ;
wire \pre_mepc[10]~q ;
wire \mepc[10]~8_combout ;
wire \_T_244[10]~12_combout ;
wire \_T_244[10]~13_combout ;
wire \pre_mepc~12_combout ;
wire \pre_mepc[11]~q ;
wire \mepc[11]~9_combout ;
wire \_T_244[11]~14_combout ;
wire \_T_244[11]~15_combout ;
wire \pre_mepc~13_combout ;
wire \pre_mepc[12]~q ;
wire \mepc[12]~10_combout ;
wire \_T_244[12]~16_combout ;
wire \_T_244[12]~17_combout ;
wire \pre_mepc~14_combout ;
wire \pre_mepc[13]~q ;
wire \mepc[13]~11_combout ;
wire \_T_244[13]~18_combout ;
wire \_T_244[13]~19_combout ;
wire \pre_mepc~15_combout ;
wire \pre_mepc[14]~q ;
wire \mepc[14]~12_combout ;
wire \_T_244[14]~20_combout ;
wire \_T_244[14]~21_combout ;
wire \pre_mepc~16_combout ;
wire \pre_mepc[15]~q ;
wire \mepc[15]~13_combout ;
wire \_T_244[15]~22_combout ;
wire \_T_244[15]~23_combout ;
wire \pre_mepc~17_combout ;
wire \pre_mepc[16]~q ;
wire \mepc[16]~14_combout ;
wire \_T_244[16]~24_combout ;
wire \_T_244[16]~25_combout ;
wire \pre_mepc~18_combout ;
wire \pre_mepc[17]~q ;
wire \mepc[17]~15_combout ;
wire \_T_244[17]~26_combout ;
wire \_T_244[17]~27_combout ;
wire \pre_mepc~19_combout ;
wire \pre_mepc[18]~q ;
wire \mepc[18]~16_combout ;
wire \_T_244[18]~28_combout ;
wire \_T_244[18]~29_combout ;
wire \pre_mepc~20_combout ;
wire \pre_mepc[19]~q ;
wire \mepc[19]~17_combout ;
wire \_T_244[19]~30_combout ;
wire \_T_244[19]~31_combout ;
wire \pre_mepc~21_combout ;
wire \pre_mepc[20]~q ;
wire \mepc[20]~18_combout ;
wire \_T_244[20]~32_combout ;
wire \_T_244[20]~33_combout ;
wire \pre_mepc~22_combout ;
wire \pre_mepc[21]~q ;
wire \mepc[21]~19_combout ;
wire \io_out[21]~195_combout ;
wire \_T_244[21]~34_combout ;
wire \_T_244[21]~35_combout ;
wire \pre_mepc~23_combout ;
wire \pre_mepc[22]~q ;
wire \mepc[22]~20_combout ;
wire \_T_244[22]~36_combout ;
wire \_T_244[22]~37_combout ;
wire \pre_mepc~24_combout ;
wire \pre_mepc[23]~q ;
wire \mepc[23]~21_combout ;
wire \_T_244[23]~38_combout ;
wire \_T_244[23]~39_combout ;
wire \pre_mepc~25_combout ;
wire \pre_mepc[24]~q ;
wire \mepc[24]~22_combout ;
wire \_T_244[24]~40_combout ;
wire \_T_244[24]~41_combout ;
wire \pre_mepc~26_combout ;
wire \pre_mepc[25]~q ;
wire \mepc[25]~23_combout ;
wire \io_out[25]~223_combout ;
wire \_T_244[25]~42_combout ;
wire \_T_244[25]~43_combout ;
wire \pre_mepc~27_combout ;
wire \pre_mepc[26]~q ;
wire \mepc[26]~24_combout ;
wire \_T_244[26]~44_combout ;
wire \_T_244[26]~45_combout ;
wire \pre_mepc~28_combout ;
wire \pre_mepc[27]~q ;
wire \mepc[27]~25_combout ;
wire \io_out[27]~237_combout ;
wire \_T_244[27]~46_combout ;
wire \_T_244[27]~47_combout ;
wire \pre_mepc~29_combout ;
wire \pre_mepc[28]~q ;
wire \mepc[28]~26_combout ;
wire \_T_244[28]~48_combout ;
wire \_T_244[28]~49_combout ;
wire \pre_mepc~30_combout ;
wire \pre_mepc[29]~q ;
wire \mepc[29]~27_combout ;
wire \io_out[29]~38_combout ;
wire \_T_244[29]~50_combout ;
wire \_T_244[29]~51_combout ;
wire \pre_mepc~31_combout ;
wire \pre_mepc[30]~q ;
wire \mepc[30]~28_combout ;
wire \_T_244[30]~52_combout ;
wire \_T_244[30]~53_combout ;
wire \pre_mepc~32_combout ;
wire \pre_mepc[31]~q ;
wire \mepc[31]~29_combout ;
wire \_T_246[31]~9_combout ;
wire \_T_246[31]~10_combout ;
wire \isIllegal~0_combout ;
wire \iaddrInvalid_j~0_combout ;
wire \mcause~4_combout ;
wire \laddrInvalid~0_combout ;
wire \saddrInvalid~0_combout ;
wire \Add0~0_combout ;
wire \Add0~1_combout ;
wire \laddrInvalid~1_combout ;
wire \mcause[0]~5_combout ;
wire \pre_mepc~0_combout ;
wire \pre_mepc[0]~q ;
wire \_GEN_204[0]~0_combout ;
wire \_T_246[0]~1_combout ;
wire \_T_246[0]~2_combout ;
wire \mtvec~0_combout ;
wire \Equal19~1_combout ;
wire \Equal19~2_combout ;
wire \Equal19~3_combout ;
wire \instreth~32_combout ;
wire \mtvec[5]~1_combout ;
wire \pre_mepc~2_combout ;
wire \pre_mepc[1]~q ;
wire \_GEN_204[1]~1_combout ;
wire \_T_246[1]~3_combout ;
wire \_T_246[1]~4_combout ;
wire \mtvec~2_combout ;
wire \Equal30~0_combout ;
wire \Equal25~3_combout ;
wire \mscratch[0]~0_combout ;
wire \mscratch[1]~q ;
wire \io_out[1]~2_combout ;
wire \Equal16~1_combout ;
wire \Equal3~0_combout ;
wire \Equal11~2_combout ;
wire \Equal11~3_combout ;
wire \Equal23~0_combout ;
wire \io_out[1]~3_combout ;
wire \io_out[1]~4_combout ;
wire \time_[0]~32_combout ;
wire \Equal19~4_combout ;
wire \Equal21~2_combout ;
wire \Equal29~2_combout ;
wire \timeh~33_combout ;
wire \time_~36_combout ;
wire \time_[0]~q ;
wire \time_[0]~33 ;
wire \time_[1]~34_combout ;
wire \time_[1]~q ;
wire \io_out[1]~5_combout ;
wire \Equal9~0_combout ;
wire \io_out[1]~6_combout ;
wire \cycle[0]~32_combout ;
wire \cycle~36_combout ;
wire \cycle[0]~q ;
wire \cycle[0]~33 ;
wire \cycle[1]~34_combout ;
wire \cycle[1]~q ;
wire \io_out[1]~7_combout ;
wire \Equal25~5_combout ;
wire \Equal27~0_combout ;
wire \Equal12~0_combout ;
wire \Equal8~0_combout ;
wire \io_out[1]~8_combout ;
wire \instret[0]~34_combout ;
wire \instret~38_combout ;
wire \Equal39~0_combout ;
wire \Equal39~1_combout ;
wire \Equal39~2_combout ;
wire \Equal39~3_combout ;
wire \Equal39~4_combout ;
wire \Equal39~5_combout ;
wire \Equal39~6_combout ;
wire \isInstRet~0_combout ;
wire \instret[0]~99_combout ;
wire \instret[0]~q ;
wire \instret[0]~35 ;
wire \instret[1]~36_combout ;
wire \instret[1]~q ;
wire \mcause[2]~7_combout ;
wire \_T_219~0_combout ;
wire \mcause~8_combout ;
wire \saddrInvalid~1_combout ;
wire \mcause~9_combout ;
wire \mcause~10_combout ;
wire \mcause[0]~11_combout ;
wire \mcause[1]~q ;
wire \io_out[1]~9_combout ;
wire \Equal28~0_combout ;
wire \Equal13~0_combout ;
wire \io_out[1]~10_combout ;
wire \cycleh[0]~32_combout ;
wire \cycleh~36_combout ;
wire \cycle[1]~35 ;
wire \cycle[2]~37_combout ;
wire \cycle[2]~q ;
wire \cycle[2]~38 ;
wire \cycle[3]~39_combout ;
wire \cycle[3]~q ;
wire \cycle[3]~40 ;
wire \cycle[4]~41_combout ;
wire \cycle[4]~q ;
wire \cycle[4]~42 ;
wire \cycle[5]~43_combout ;
wire \cycle[5]~q ;
wire \cycle[5]~44 ;
wire \cycle[6]~45_combout ;
wire \cycle[6]~q ;
wire \cycle[6]~46 ;
wire \cycle[7]~47_combout ;
wire \cycle[7]~q ;
wire \cycle[7]~48 ;
wire \cycle[8]~49_combout ;
wire \cycle[8]~q ;
wire \cycle[8]~50 ;
wire \cycle[9]~51_combout ;
wire \cycle[9]~q ;
wire \cycle[9]~52 ;
wire \cycle[10]~53_combout ;
wire \cycle[10]~q ;
wire \cycle[10]~54 ;
wire \cycle[11]~55_combout ;
wire \cycle[11]~q ;
wire \cycle[11]~56 ;
wire \cycle[12]~57_combout ;
wire \cycle[12]~q ;
wire \cycle[12]~58 ;
wire \cycle[13]~59_combout ;
wire \cycle[13]~q ;
wire \cycle[13]~60 ;
wire \cycle[14]~61_combout ;
wire \cycle[14]~q ;
wire \cycle[14]~62 ;
wire \cycle[15]~63_combout ;
wire \cycle[15]~q ;
wire \cycle[15]~64 ;
wire \cycle[16]~65_combout ;
wire \cycle[16]~q ;
wire \cycle[16]~66 ;
wire \cycle[17]~67_combout ;
wire \cycle[17]~q ;
wire \cycle[17]~68 ;
wire \cycle[18]~69_combout ;
wire \cycle[18]~q ;
wire \cycle[18]~70 ;
wire \cycle[19]~71_combout ;
wire \cycle[19]~q ;
wire \cycle[19]~72 ;
wire \cycle[20]~73_combout ;
wire \cycle[20]~q ;
wire \cycle[20]~74 ;
wire \cycle[21]~75_combout ;
wire \cycle[21]~q ;
wire \cycle[21]~76 ;
wire \cycle[22]~77_combout ;
wire \cycle[22]~q ;
wire \cycle[22]~78 ;
wire \cycle[23]~79_combout ;
wire \cycle[23]~q ;
wire \cycle[23]~80 ;
wire \cycle[24]~81_combout ;
wire \cycle[24]~q ;
wire \cycle[24]~82 ;
wire \cycle[25]~83_combout ;
wire \cycle[25]~q ;
wire \cycle[25]~84 ;
wire \cycle[26]~85_combout ;
wire \cycle[26]~q ;
wire \cycle[26]~86 ;
wire \cycle[27]~87_combout ;
wire \cycle[27]~q ;
wire \cycle[27]~88 ;
wire \cycle[28]~89_combout ;
wire \cycle[28]~q ;
wire \cycle[28]~90 ;
wire \cycle[29]~91_combout ;
wire \cycle[29]~q ;
wire \cycle[29]~92 ;
wire \cycle[30]~93_combout ;
wire \cycle[30]~q ;
wire \cycle[30]~94 ;
wire \cycle[31]~95_combout ;
wire \cycle[31]~q ;
wire \WideAnd1~0_combout ;
wire \WideAnd1~1_combout ;
wire \WideAnd1~2_combout ;
wire \WideAnd1~3_combout ;
wire \WideAnd1~4_combout ;
wire \WideAnd1~5_combout ;
wire \WideAnd1~6_combout ;
wire \WideAnd1~7_combout ;
wire \WideAnd1~8_combout ;
wire \WideAnd1~9_combout ;
wire \cycleh[23]~37_combout ;
wire \cycleh[0]~q ;
wire \cycleh[0]~33 ;
wire \cycleh[1]~34_combout ;
wire \cycleh[1]~q ;
wire \mbadaddr[0]~0_combout ;
wire \mbadaddr[1]~q ;
wire \io_out[1]~11_combout ;
wire \timeh~32_combout ;
wire \io_out[1]~12_combout ;
wire \timeh[0]~34_combout ;
wire \timeh~38_combout ;
wire \time_[1]~35 ;
wire \time_[2]~37_combout ;
wire \time_[2]~q ;
wire \time_[2]~38 ;
wire \time_[3]~39_combout ;
wire \time_[3]~q ;
wire \time_[3]~40 ;
wire \time_[4]~41_combout ;
wire \time_[4]~q ;
wire \time_[4]~42 ;
wire \time_[5]~43_combout ;
wire \time_[5]~q ;
wire \time_[5]~44 ;
wire \time_[6]~45_combout ;
wire \time_[6]~q ;
wire \time_[6]~46 ;
wire \time_[7]~47_combout ;
wire \time_[7]~q ;
wire \time_[7]~48 ;
wire \time_[8]~49_combout ;
wire \time_[8]~q ;
wire \time_[8]~50 ;
wire \time_[9]~51_combout ;
wire \time_[9]~q ;
wire \time_[9]~52 ;
wire \time_[10]~53_combout ;
wire \time_[10]~q ;
wire \time_[10]~54 ;
wire \time_[11]~55_combout ;
wire \time_[11]~q ;
wire \time_[11]~56 ;
wire \time_[12]~57_combout ;
wire \time_[12]~q ;
wire \time_[12]~58 ;
wire \time_[13]~59_combout ;
wire \time_[13]~q ;
wire \time_[13]~60 ;
wire \time_[14]~61_combout ;
wire \time_[14]~q ;
wire \time_[14]~62 ;
wire \time_[15]~63_combout ;
wire \time_[15]~q ;
wire \time_[15]~64 ;
wire \time_[16]~65_combout ;
wire \time_[16]~q ;
wire \time_[16]~66 ;
wire \time_[17]~67_combout ;
wire \time_[17]~q ;
wire \time_[17]~68 ;
wire \time_[18]~69_combout ;
wire \time_[18]~q ;
wire \time_[18]~70 ;
wire \time_[19]~71_combout ;
wire \time_[19]~q ;
wire \time_[19]~72 ;
wire \time_[20]~73_combout ;
wire \time_[20]~q ;
wire \time_[20]~74 ;
wire \time_[21]~75_combout ;
wire \time_[21]~q ;
wire \time_[21]~76 ;
wire \time_[22]~77_combout ;
wire \time_[22]~q ;
wire \time_[22]~78 ;
wire \time_[23]~79_combout ;
wire \time_[23]~q ;
wire \time_[23]~80 ;
wire \time_[24]~81_combout ;
wire \time_[24]~q ;
wire \time_[24]~82 ;
wire \time_[25]~83_combout ;
wire \time_[25]~q ;
wire \time_[25]~84 ;
wire \time_[26]~85_combout ;
wire \time_[26]~q ;
wire \time_[26]~86 ;
wire \time_[27]~87_combout ;
wire \time_[27]~q ;
wire \time_[27]~88 ;
wire \time_[28]~89_combout ;
wire \time_[28]~q ;
wire \time_[28]~90 ;
wire \time_[29]~91_combout ;
wire \time_[29]~q ;
wire \time_[29]~92 ;
wire \time_[30]~93_combout ;
wire \time_[30]~q ;
wire \time_[30]~94 ;
wire \time_[31]~95_combout ;
wire \time_[31]~q ;
wire \WideAnd0~0_combout ;
wire \WideAnd0~1_combout ;
wire \WideAnd0~2_combout ;
wire \WideAnd0~3_combout ;
wire \WideAnd0~4_combout ;
wire \WideAnd0~5_combout ;
wire \WideAnd0~6_combout ;
wire \WideAnd0~7_combout ;
wire \WideAnd0~8_combout ;
wire \WideAnd0~9_combout ;
wire \timeh[31]~39_combout ;
wire \timeh[0]~q ;
wire \timeh[0]~35 ;
wire \timeh[1]~36_combout ;
wire \timeh[1]~q ;
wire \io_out[1]~13_combout ;
wire \Equal13~1_combout ;
wire \io_out[1]~14_combout ;
wire \instreth[0]~33_combout ;
wire \instreth~37_combout ;
wire \isInstRet~combout ;
wire \instret[1]~37 ;
wire \instret[2]~39_combout ;
wire \instret[2]~q ;
wire \instret[2]~40 ;
wire \instret[3]~41_combout ;
wire \instret[3]~q ;
wire \instret[3]~42 ;
wire \instret[4]~43_combout ;
wire \instret[4]~q ;
wire \instret[4]~44 ;
wire \instret[5]~45_combout ;
wire \instret[5]~q ;
wire \instret[5]~46 ;
wire \instret[6]~47_combout ;
wire \instret[6]~q ;
wire \instret[6]~48 ;
wire \instret[7]~49_combout ;
wire \instret[7]~q ;
wire \instret[7]~50 ;
wire \instret[8]~51_combout ;
wire \instret[8]~q ;
wire \instret[8]~52 ;
wire \instret[9]~53_combout ;
wire \instret[9]~q ;
wire \instret[9]~54 ;
wire \instret[10]~55_combout ;
wire \instret[10]~q ;
wire \instret[10]~56 ;
wire \instret[11]~57_combout ;
wire \instret[11]~q ;
wire \instret[11]~58 ;
wire \instret[12]~59_combout ;
wire \instret[12]~q ;
wire \instret[12]~60 ;
wire \instret[13]~61_combout ;
wire \instret[13]~q ;
wire \instret[13]~62 ;
wire \instret[14]~63_combout ;
wire \instret[14]~q ;
wire \instret[14]~64 ;
wire \instret[15]~65_combout ;
wire \instret[15]~q ;
wire \instret[15]~66 ;
wire \instret[16]~67_combout ;
wire \instret[16]~q ;
wire \instret[16]~68 ;
wire \instret[17]~69_combout ;
wire \instret[17]~q ;
wire \instret[17]~70 ;
wire \instret[18]~71_combout ;
wire \instret[18]~q ;
wire \instret[18]~72 ;
wire \instret[19]~73_combout ;
wire \instret[19]~q ;
wire \instret[19]~74 ;
wire \instret[20]~75_combout ;
wire \instret[20]~q ;
wire \instret[20]~76 ;
wire \instret[21]~77_combout ;
wire \instret[21]~q ;
wire \instret[21]~78 ;
wire \instret[22]~79_combout ;
wire \instret[22]~q ;
wire \instret[22]~80 ;
wire \instret[23]~81_combout ;
wire \instret[23]~q ;
wire \instret[23]~82 ;
wire \instret[24]~83_combout ;
wire \instret[24]~q ;
wire \instret[24]~84 ;
wire \instret[25]~85_combout ;
wire \instret[25]~q ;
wire \instret[25]~86 ;
wire \instret[26]~87_combout ;
wire \instret[26]~q ;
wire \instret[26]~88 ;
wire \instret[27]~89_combout ;
wire \instret[27]~q ;
wire \instret[27]~90 ;
wire \instret[28]~91_combout ;
wire \instret[28]~q ;
wire \instret[28]~92 ;
wire \instret[29]~93_combout ;
wire \instret[29]~q ;
wire \instret[29]~94 ;
wire \instret[30]~95_combout ;
wire \instret[30]~q ;
wire \instret[30]~96 ;
wire \instret[31]~97_combout ;
wire \instret[31]~q ;
wire \_T_198~0_combout ;
wire \_T_198~1_combout ;
wire \_T_198~2_combout ;
wire \_T_198~3_combout ;
wire \_T_198~4_combout ;
wire \_T_198~5_combout ;
wire \_T_198~6_combout ;
wire \_T_198~7_combout ;
wire \_T_198~8_combout ;
wire \_T_198~9_combout ;
wire \_T_198~combout ;
wire \instreth[3]~38_combout ;
wire \instreth[0]~q ;
wire \instreth[0]~34 ;
wire \instreth[1]~35_combout ;
wire \instreth[1]~q ;
wire \io_out[1]~15_combout ;
wire \mscratch[0]~q ;
wire \io_out[0]~17_combout ;
wire \io_out[0]~18_combout ;
wire \mcause[0]~12_combout ;
wire \mcause[0]~q ;
wire \io_out[0]~19_combout ;
wire \mbadaddr[0]~q ;
wire \io_out[0]~20_combout ;
wire \io_out[0]~21_combout ;
wire \IE~2_combout ;
wire \IE1~0_combout ;
wire \PRV1[0]~4_combout ;
wire \IE~q ;
wire \io_out[0]~22_combout ;
wire \io_out[0]~23_combout ;
wire \mtvec~3_combout ;
wire \mtvec~4_combout ;
wire \mtvec~5_combout ;
wire \mtvec~6_combout ;
wire \mtvec~7_combout ;
wire \mtvec~8_combout ;
wire \mtvec~9_combout ;
wire \mtvec~10_combout ;
wire \mtvec~11_combout ;
wire \mtvec~12_combout ;
wire \mtvec~13_combout ;
wire \mtvec~14_combout ;
wire \mtvec~15_combout ;
wire \mtvec~16_combout ;
wire \mtvec~17_combout ;
wire \mtvec~18_combout ;
wire \mtvec~19_combout ;
wire \mtvec~20_combout ;
wire \mtvec~21_combout ;
wire \mtvec~22_combout ;
wire \mtvec~23_combout ;
wire \mtvec~24_combout ;
wire \mtvec~25_combout ;
wire \mtvec~26_combout ;
wire \mtvec~27_combout ;
wire \mtvec~28_combout ;
wire \mtvec~29_combout ;
wire \mtvec~30_combout ;
wire \mtvec~31_combout ;
wire \mtvec~32_combout ;
wire \mscratch[28]~q ;
wire \io_out[28]~25_combout ;
wire \io_out[28]~26_combout ;
wire \mbadaddr[28]~q ;
wire \io_out[28]~27_combout ;
wire \cycleh[1]~35 ;
wire \cycleh[2]~38_combout ;
wire \cycleh[2]~q ;
wire \cycleh[2]~39 ;
wire \cycleh[3]~40_combout ;
wire \cycleh[3]~q ;
wire \cycleh[3]~41 ;
wire \cycleh[4]~42_combout ;
wire \cycleh[4]~q ;
wire \cycleh[4]~43 ;
wire \cycleh[5]~44_combout ;
wire \cycleh[5]~q ;
wire \cycleh[5]~45 ;
wire \cycleh[6]~46_combout ;
wire \cycleh[6]~q ;
wire \cycleh[6]~47 ;
wire \cycleh[7]~48_combout ;
wire \cycleh[7]~q ;
wire \cycleh[7]~49 ;
wire \cycleh[8]~50_combout ;
wire \cycleh[8]~q ;
wire \cycleh[8]~51 ;
wire \cycleh[9]~52_combout ;
wire \cycleh[9]~q ;
wire \cycleh[9]~53 ;
wire \cycleh[10]~54_combout ;
wire \cycleh[10]~q ;
wire \cycleh[10]~55 ;
wire \cycleh[11]~56_combout ;
wire \cycleh[11]~q ;
wire \cycleh[11]~57 ;
wire \cycleh[12]~58_combout ;
wire \cycleh[12]~q ;
wire \cycleh[12]~59 ;
wire \cycleh[13]~60_combout ;
wire \cycleh[13]~q ;
wire \cycleh[13]~61 ;
wire \cycleh[14]~62_combout ;
wire \cycleh[14]~q ;
wire \cycleh[14]~63 ;
wire \cycleh[15]~64_combout ;
wire \cycleh[15]~q ;
wire \cycleh[15]~65 ;
wire \cycleh[16]~66_combout ;
wire \cycleh[16]~q ;
wire \cycleh[16]~67 ;
wire \cycleh[17]~68_combout ;
wire \cycleh[17]~q ;
wire \cycleh[17]~69 ;
wire \cycleh[18]~70_combout ;
wire \cycleh[18]~q ;
wire \cycleh[18]~71 ;
wire \cycleh[19]~72_combout ;
wire \cycleh[19]~q ;
wire \cycleh[19]~73 ;
wire \cycleh[20]~74_combout ;
wire \cycleh[20]~q ;
wire \cycleh[20]~75 ;
wire \cycleh[21]~76_combout ;
wire \cycleh[21]~q ;
wire \cycleh[21]~77 ;
wire \cycleh[22]~78_combout ;
wire \cycleh[22]~q ;
wire \cycleh[22]~79 ;
wire \cycleh[23]~80_combout ;
wire \cycleh[23]~q ;
wire \cycleh[23]~81 ;
wire \cycleh[24]~82_combout ;
wire \cycleh[24]~q ;
wire \cycleh[24]~83 ;
wire \cycleh[25]~84_combout ;
wire \cycleh[25]~q ;
wire \cycleh[25]~85 ;
wire \cycleh[26]~86_combout ;
wire \cycleh[26]~q ;
wire \cycleh[26]~87 ;
wire \cycleh[27]~88_combout ;
wire \cycleh[27]~q ;
wire \cycleh[27]~89 ;
wire \cycleh[28]~90_combout ;
wire \cycleh[28]~q ;
wire \io_out[28]~28_combout ;
wire \io_out[28]~29_combout ;
wire \instreth[1]~36 ;
wire \instreth[2]~39_combout ;
wire \instreth[2]~q ;
wire \instreth[2]~40 ;
wire \instreth[3]~41_combout ;
wire \instreth[3]~q ;
wire \instreth[3]~42 ;
wire \instreth[4]~43_combout ;
wire \instreth[4]~q ;
wire \instreth[4]~44 ;
wire \instreth[5]~45_combout ;
wire \instreth[5]~q ;
wire \instreth[5]~46 ;
wire \instreth[6]~47_combout ;
wire \instreth[6]~q ;
wire \instreth[6]~48 ;
wire \instreth[7]~49_combout ;
wire \instreth[7]~q ;
wire \instreth[7]~50 ;
wire \instreth[8]~51_combout ;
wire \instreth[8]~q ;
wire \instreth[8]~52 ;
wire \instreth[9]~53_combout ;
wire \instreth[9]~q ;
wire \instreth[9]~54 ;
wire \instreth[10]~55_combout ;
wire \instreth[10]~q ;
wire \instreth[10]~56 ;
wire \instreth[11]~57_combout ;
wire \instreth[11]~q ;
wire \instreth[11]~58 ;
wire \instreth[12]~59_combout ;
wire \instreth[12]~q ;
wire \instreth[12]~60 ;
wire \instreth[13]~61_combout ;
wire \instreth[13]~q ;
wire \instreth[13]~62 ;
wire \instreth[14]~63_combout ;
wire \instreth[14]~q ;
wire \instreth[14]~64 ;
wire \instreth[15]~65_combout ;
wire \instreth[15]~q ;
wire \instreth[15]~66 ;
wire \instreth[16]~67_combout ;
wire \instreth[16]~q ;
wire \instreth[16]~68 ;
wire \instreth[17]~69_combout ;
wire \instreth[17]~q ;
wire \instreth[17]~70 ;
wire \instreth[18]~71_combout ;
wire \instreth[18]~q ;
wire \instreth[18]~72 ;
wire \instreth[19]~73_combout ;
wire \instreth[19]~q ;
wire \instreth[19]~74 ;
wire \instreth[20]~75_combout ;
wire \instreth[20]~q ;
wire \instreth[20]~76 ;
wire \instreth[21]~77_combout ;
wire \instreth[21]~q ;
wire \instreth[21]~78 ;
wire \instreth[22]~79_combout ;
wire \instreth[22]~q ;
wire \instreth[22]~80 ;
wire \instreth[23]~81_combout ;
wire \instreth[23]~q ;
wire \instreth[23]~82 ;
wire \instreth[24]~83_combout ;
wire \instreth[24]~q ;
wire \instreth[24]~84 ;
wire \instreth[25]~85_combout ;
wire \instreth[25]~q ;
wire \instreth[25]~86 ;
wire \instreth[26]~87_combout ;
wire \instreth[26]~q ;
wire \instreth[26]~88 ;
wire \instreth[27]~89_combout ;
wire \instreth[27]~q ;
wire \instreth[27]~90 ;
wire \instreth[28]~91_combout ;
wire \instreth[28]~q ;
wire \io_out[28]~30_combout ;
wire \timeh[1]~37 ;
wire \timeh[2]~40_combout ;
wire \timeh[2]~q ;
wire \timeh[2]~41 ;
wire \timeh[3]~42_combout ;
wire \timeh[3]~q ;
wire \timeh[3]~43 ;
wire \timeh[4]~44_combout ;
wire \timeh[4]~q ;
wire \timeh[4]~45 ;
wire \timeh[5]~46_combout ;
wire \timeh[5]~q ;
wire \timeh[5]~47 ;
wire \timeh[6]~48_combout ;
wire \timeh[6]~q ;
wire \timeh[6]~49 ;
wire \timeh[7]~50_combout ;
wire \timeh[7]~q ;
wire \timeh[7]~51 ;
wire \timeh[8]~52_combout ;
wire \timeh[8]~q ;
wire \timeh[8]~53 ;
wire \timeh[9]~54_combout ;
wire \timeh[9]~q ;
wire \timeh[9]~55 ;
wire \timeh[10]~56_combout ;
wire \timeh[10]~q ;
wire \timeh[10]~57 ;
wire \timeh[11]~58_combout ;
wire \timeh[11]~q ;
wire \timeh[11]~59 ;
wire \timeh[12]~60_combout ;
wire \timeh[12]~q ;
wire \timeh[12]~61 ;
wire \timeh[13]~62_combout ;
wire \timeh[13]~q ;
wire \timeh[13]~63 ;
wire \timeh[14]~64_combout ;
wire \timeh[14]~q ;
wire \timeh[14]~65 ;
wire \timeh[15]~66_combout ;
wire \timeh[15]~q ;
wire \timeh[15]~67 ;
wire \timeh[16]~68_combout ;
wire \timeh[16]~q ;
wire \timeh[16]~69 ;
wire \timeh[17]~70_combout ;
wire \timeh[17]~q ;
wire \timeh[17]~71 ;
wire \timeh[18]~72_combout ;
wire \timeh[18]~q ;
wire \timeh[18]~73 ;
wire \timeh[19]~74_combout ;
wire \timeh[19]~q ;
wire \timeh[19]~75 ;
wire \timeh[20]~76_combout ;
wire \timeh[20]~q ;
wire \timeh[20]~77 ;
wire \timeh[21]~78_combout ;
wire \timeh[21]~q ;
wire \timeh[21]~79 ;
wire \timeh[22]~80_combout ;
wire \timeh[22]~q ;
wire \timeh[22]~81 ;
wire \timeh[23]~82_combout ;
wire \timeh[23]~q ;
wire \timeh[23]~83 ;
wire \timeh[24]~84_combout ;
wire \timeh[24]~q ;
wire \timeh[24]~85 ;
wire \timeh[25]~86_combout ;
wire \timeh[25]~q ;
wire \timeh[25]~87 ;
wire \timeh[26]~88_combout ;
wire \timeh[26]~q ;
wire \timeh[26]~89 ;
wire \timeh[27]~90_combout ;
wire \timeh[27]~q ;
wire \timeh[27]~91 ;
wire \timeh[28]~92_combout ;
wire \timeh[28]~q ;
wire \mscratch[29]~q ;
wire \io_out[29]~32_combout ;
wire \io_out[29]~33_combout ;
wire \mbadaddr[29]~q ;
wire \io_out[29]~34_combout ;
wire \cycleh[28]~91 ;
wire \cycleh[29]~92_combout ;
wire \cycleh[29]~q ;
wire \io_out[29]~35_combout ;
wire \instreth[28]~92 ;
wire \instreth[29]~93_combout ;
wire \instreth[29]~q ;
wire \timeh[28]~93 ;
wire \timeh[29]~94_combout ;
wire \timeh[29]~q ;
wire \mscratch[30]~q ;
wire \io_out[30]~39_combout ;
wire \io_out[30]~40_combout ;
wire \io_out[30]~41_combout ;
wire \mbadaddr[30]~q ;
wire \io_out[30]~42_combout ;
wire \cycleh[29]~93 ;
wire \cycleh[30]~94_combout ;
wire \cycleh[30]~q ;
wire \io_out[30]~43_combout ;
wire \instreth[29]~94 ;
wire \instreth[30]~95_combout ;
wire \instreth[30]~q ;
wire \timeh[29]~95 ;
wire \timeh[30]~96_combout ;
wire \timeh[30]~q ;
wire \io_out[30]~44_combout ;
wire \mscratch[31]~q ;
wire \io_out[31]~46_combout ;
wire \io_out[31]~47_combout ;
wire \mcause[31]~13_combout ;
wire \mcause[31]~q ;
wire \io_out[31]~48_combout ;
wire \cycleh[30]~95 ;
wire \cycleh[31]~96_combout ;
wire \cycleh[31]~q ;
wire \mbadaddr[31]~q ;
wire \io_out[31]~49_combout ;
wire \io_out[31]~50_combout ;
wire \timeh[30]~97 ;
wire \timeh[31]~98_combout ;
wire \timeh[31]~q ;
wire \io_out[31]~51_combout ;
wire \instreth[30]~96 ;
wire \instreth[31]~97_combout ;
wire \instreth[31]~q ;
wire \Equal16~2_combout ;
wire \mscratch[8]~q ;
wire \io_out[8]~53_combout ;
wire \io_out[8]~54_combout ;
wire \io_out[8]~55_combout ;
wire \mbadaddr[8]~q ;
wire \io_out[8]~56_combout ;
wire \io_out[8]~57_combout ;
wire \io_out[8]~58_combout ;
wire \mscratch[9]~q ;
wire \io_out[9]~60_combout ;
wire \io_out[9]~61_combout ;
wire \mbadaddr[9]~q ;
wire \io_out[9]~62_combout ;
wire \io_out[9]~63_combout ;
wire \io_out[9]~64_combout ;
wire \io_out[9]~65_combout ;
wire \mscratch[10]~q ;
wire \io_out[10]~67_combout ;
wire \Equal25~4_combout ;
wire \io_out[10]~238_combout ;
wire \io_out[10]~68_combout ;
wire \mbadaddr[10]~q ;
wire \io_out[10]~69_combout ;
wire \io_out[10]~70_combout ;
wire \io_out[10]~71_combout ;
wire \mscratch[11]~q ;
wire \io_out[11]~73_combout ;
wire \io_out[11]~74_combout ;
wire \mbadaddr[11]~q ;
wire \io_out[11]~75_combout ;
wire \MTIE~0_combout ;
wire \MEIE~q ;
wire \io_out[11]~76_combout ;
wire \io_out[11]~77_combout ;
wire \io_out[11]~78_combout ;
wire \mscratch[12]~q ;
wire \io_out[12]~80_combout ;
wire \io_out[12]~81_combout ;
wire \io_out[12]~82_combout ;
wire \mbadaddr[12]~q ;
wire \io_out[12]~83_combout ;
wire \io_out[12]~84_combout ;
wire \io_out[12]~85_combout ;
wire \mscratch[13]~q ;
wire \io_out[13]~87_combout ;
wire \io_out[13]~88_combout ;
wire \mbadaddr[13]~q ;
wire \io_out[13]~89_combout ;
wire \io_out[13]~90_combout ;
wire \io_out[13]~91_combout ;
wire \io_out[13]~92_combout ;
wire \mscratch[14]~q ;
wire \io_out[14]~94_combout ;
wire \io_out[14]~95_combout ;
wire \io_out[14]~96_combout ;
wire \mbadaddr[14]~q ;
wire \io_out[14]~97_combout ;
wire \io_out[14]~98_combout ;
wire \io_out[14]~99_combout ;
wire \mscratch[15]~q ;
wire \io_out[15]~101_combout ;
wire \io_out[15]~102_combout ;
wire \mbadaddr[15]~q ;
wire \io_out[15]~103_combout ;
wire \io_out[15]~104_combout ;
wire \io_out[15]~105_combout ;
wire \io_out[15]~106_combout ;
wire \mscratch[16]~q ;
wire \io_out[16]~108_combout ;
wire \io_out[16]~109_combout ;
wire \io_out[16]~110_combout ;
wire \mbadaddr[16]~q ;
wire \io_out[16]~111_combout ;
wire \io_out[16]~112_combout ;
wire \io_out[16]~113_combout ;
wire \mscratch[17]~q ;
wire \io_out[17]~115_combout ;
wire \io_out[17]~116_combout ;
wire \io_out[17]~117_combout ;
wire \mbadaddr[17]~q ;
wire \io_out[17]~118_combout ;
wire \io_out[17]~119_combout ;
wire \io_out[17]~120_combout ;
wire \mscratch[18]~q ;
wire \io_out[18]~122_combout ;
wire \io_out[18]~123_combout ;
wire \mbadaddr[18]~q ;
wire \io_out[18]~124_combout ;
wire \io_out[18]~125_combout ;
wire \io_out[18]~126_combout ;
wire \io_out[18]~127_combout ;
wire \mscratch[19]~q ;
wire \io_out[19]~129_combout ;
wire \io_out[19]~130_combout ;
wire \mbadaddr[19]~q ;
wire \io_out[19]~131_combout ;
wire \io_out[19]~132_combout ;
wire \io_out[19]~133_combout ;
wire \io_out[19]~134_combout ;
wire \mscratch[4]~q ;
wire \io_out[4]~136_combout ;
wire \io_out[4]~137_combout ;
wire \mbadaddr[4]~q ;
wire \io_out[4]~138_combout ;
wire \PRV1~5_combout ;
wire \PRV1[0]~q ;
wire \io_out[4]~139_combout ;
wire \io_out[4]~140_combout ;
wire \io_out[4]~141_combout ;
wire \mscratch[2]~q ;
wire \io_out[2]~143_combout ;
wire \io_out[2]~144_combout ;
wire \io_out[2]~145_combout ;
wire \mcause~14_combout ;
wire \mcause~15_combout ;
wire \mcause[2]~q ;
wire \io_out[2]~146_combout ;
wire \mbadaddr[2]~q ;
wire \io_out[2]~147_combout ;
wire \io_out[2]~148_combout ;
wire \io_out[2]~149_combout ;
wire \MSIE~q ;
wire \io_out[3]~151_combout ;
wire \mscratch[3]~q ;
wire \io_out[3]~152_combout ;
wire \io_out[3]~153_combout ;
wire \io_out[3]~154_combout ;
wire \mcause[3]~16_combout ;
wire \mcause[3]~q ;
wire \io_out[3]~155_combout ;
wire \mbadaddr[3]~q ;
wire \io_out[3]~156_combout ;
wire \MTIP~0_combout ;
wire \MSIP~q ;
wire \IE1~1_combout ;
wire \IE1~2_combout ;
wire \IE1~3_combout ;
wire \IE1~q ;
wire \io_out[3]~157_combout ;
wire \io_out[3]~158_combout ;
wire \mscratch[5]~q ;
wire \io_out[5]~160_combout ;
wire \io_out[5]~161_combout ;
wire \mbadaddr[5]~q ;
wire \io_out[5]~162_combout ;
wire \PRV1~6_combout ;
wire \PRV1[1]~q ;
wire \io_out[5]~163_combout ;
wire \io_out[5]~164_combout ;
wire \io_out[5]~165_combout ;
wire \mscratch[6]~q ;
wire \io_out[6]~167_combout ;
wire \io_out[6]~168_combout ;
wire \mbadaddr[6]~q ;
wire \io_out[6]~169_combout ;
wire \io_out[6]~170_combout ;
wire \io_out[6]~171_combout ;
wire \io_out[6]~172_combout ;
wire \MTIE~1_combout ;
wire \MTIE~q ;
wire \io_out[7]~174_combout ;
wire \io_out[7]~175_combout ;
wire \mscratch[7]~q ;
wire \io_out[7]~176_combout ;
wire \io_out[7]~177_combout ;
wire \mbadaddr[7]~q ;
wire \io_out[7]~178_combout ;
wire \io_out[7]~179_combout ;
wire \MTIP~q ;
wire \io_out[7]~180_combout ;
wire \mscratch[20]~q ;
wire \io_out[20]~182_combout ;
wire \io_out[20]~183_combout ;
wire \io_out[20]~184_combout ;
wire \mbadaddr[20]~q ;
wire \io_out[20]~185_combout ;
wire \io_out[20]~186_combout ;
wire \io_out[20]~187_combout ;
wire \mscratch[21]~q ;
wire \io_out[21]~189_combout ;
wire \io_out[21]~190_combout ;
wire \mbadaddr[21]~q ;
wire \io_out[21]~191_combout ;
wire \io_out[21]~192_combout ;
wire \mscratch[22]~q ;
wire \io_out[22]~196_combout ;
wire \io_out[22]~197_combout ;
wire \mbadaddr[22]~q ;
wire \io_out[22]~198_combout ;
wire \io_out[22]~199_combout ;
wire \io_out[22]~200_combout ;
wire \io_out[22]~201_combout ;
wire \mscratch[23]~q ;
wire \io_out[23]~203_combout ;
wire \io_out[23]~204_combout ;
wire \io_out[23]~205_combout ;
wire \mbadaddr[23]~q ;
wire \io_out[23]~206_combout ;
wire \io_out[23]~207_combout ;
wire \io_out[23]~208_combout ;
wire \mscratch[24]~q ;
wire \io_out[24]~210_combout ;
wire \io_out[24]~211_combout ;
wire \mbadaddr[24]~q ;
wire \io_out[24]~212_combout ;
wire \io_out[24]~213_combout ;
wire \io_out[24]~214_combout ;
wire \io_out[24]~215_combout ;
wire \mscratch[25]~q ;
wire \io_out[25]~217_combout ;
wire \io_out[25]~218_combout ;
wire \mbadaddr[25]~q ;
wire \io_out[25]~219_combout ;
wire \io_out[25]~220_combout ;
wire \mscratch[26]~q ;
wire \io_out[26]~224_combout ;
wire \io_out[26]~225_combout ;
wire \io_out[26]~226_combout ;
wire \mbadaddr[26]~q ;
wire \io_out[26]~227_combout ;
wire \io_out[26]~228_combout ;
wire \io_out[26]~229_combout ;
wire \mscratch[27]~q ;
wire \io_out[27]~231_combout ;
wire \io_out[27]~232_combout ;
wire \mbadaddr[27]~q ;
wire \io_out[27]~233_combout ;
wire \io_out[27]~234_combout ;


dffeas \mepc[2] (
	.clk(clock),
	.d(\mepc[2]~0_combout ),
	.asdata(\_T_246[2]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_2),
	.prn(vcc));
defparam \mepc[2] .is_wysiwyg = "true";
defparam \mepc[2] .power_up = "low";

dffeas \mepc[3] (
	.clk(clock),
	.d(\mepc[3]~1_combout ),
	.asdata(\_T_246[3]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_3),
	.prn(vcc));
defparam \mepc[3] .is_wysiwyg = "true";
defparam \mepc[3] .power_up = "low";

dffeas \mepc[4] (
	.clk(clock),
	.d(\mepc[4]~2_combout ),
	.asdata(\_T_244[4]~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_4),
	.prn(vcc));
defparam \mepc[4] .is_wysiwyg = "true";
defparam \mepc[4] .power_up = "low";

dffeas \mepc[5] (
	.clk(clock),
	.d(\mepc[5]~3_combout ),
	.asdata(\_T_244[5]~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_5),
	.prn(vcc));
defparam \mepc[5] .is_wysiwyg = "true";
defparam \mepc[5] .power_up = "low";

dffeas \mepc[6] (
	.clk(clock),
	.d(\mepc[6]~4_combout ),
	.asdata(\_T_244[6]~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_6),
	.prn(vcc));
defparam \mepc[6] .is_wysiwyg = "true";
defparam \mepc[6] .power_up = "low";

dffeas \mepc[7] (
	.clk(clock),
	.d(\mepc[7]~5_combout ),
	.asdata(\_T_244[7]~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_7),
	.prn(vcc));
defparam \mepc[7] .is_wysiwyg = "true";
defparam \mepc[7] .power_up = "low";

dffeas \mepc[8] (
	.clk(clock),
	.d(\mepc[8]~6_combout ),
	.asdata(\_T_244[8]~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_8),
	.prn(vcc));
defparam \mepc[8] .is_wysiwyg = "true";
defparam \mepc[8] .power_up = "low";

dffeas \mepc[9] (
	.clk(clock),
	.d(\mepc[9]~7_combout ),
	.asdata(\_T_244[9]~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_9),
	.prn(vcc));
defparam \mepc[9] .is_wysiwyg = "true";
defparam \mepc[9] .power_up = "low";

dffeas \mepc[10] (
	.clk(clock),
	.d(\mepc[10]~8_combout ),
	.asdata(\_T_244[10]~13_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_10),
	.prn(vcc));
defparam \mepc[10] .is_wysiwyg = "true";
defparam \mepc[10] .power_up = "low";

dffeas \mepc[11] (
	.clk(clock),
	.d(\mepc[11]~9_combout ),
	.asdata(\_T_244[11]~15_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_11),
	.prn(vcc));
defparam \mepc[11] .is_wysiwyg = "true";
defparam \mepc[11] .power_up = "low";

dffeas \mepc[12] (
	.clk(clock),
	.d(\mepc[12]~10_combout ),
	.asdata(\_T_244[12]~17_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_12),
	.prn(vcc));
defparam \mepc[12] .is_wysiwyg = "true";
defparam \mepc[12] .power_up = "low";

dffeas \mepc[13] (
	.clk(clock),
	.d(\mepc[13]~11_combout ),
	.asdata(\_T_244[13]~19_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_13),
	.prn(vcc));
defparam \mepc[13] .is_wysiwyg = "true";
defparam \mepc[13] .power_up = "low";

dffeas \mepc[14] (
	.clk(clock),
	.d(\mepc[14]~12_combout ),
	.asdata(\_T_244[14]~21_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_14),
	.prn(vcc));
defparam \mepc[14] .is_wysiwyg = "true";
defparam \mepc[14] .power_up = "low";

dffeas \mepc[15] (
	.clk(clock),
	.d(\mepc[15]~13_combout ),
	.asdata(\_T_244[15]~23_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_15),
	.prn(vcc));
defparam \mepc[15] .is_wysiwyg = "true";
defparam \mepc[15] .power_up = "low";

dffeas \mepc[16] (
	.clk(clock),
	.d(\mepc[16]~14_combout ),
	.asdata(\_T_244[16]~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_16),
	.prn(vcc));
defparam \mepc[16] .is_wysiwyg = "true";
defparam \mepc[16] .power_up = "low";

dffeas \mepc[17] (
	.clk(clock),
	.d(\mepc[17]~15_combout ),
	.asdata(\_T_244[17]~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_17),
	.prn(vcc));
defparam \mepc[17] .is_wysiwyg = "true";
defparam \mepc[17] .power_up = "low";

dffeas \mepc[18] (
	.clk(clock),
	.d(\mepc[18]~16_combout ),
	.asdata(\_T_244[18]~29_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_18),
	.prn(vcc));
defparam \mepc[18] .is_wysiwyg = "true";
defparam \mepc[18] .power_up = "low";

dffeas \mepc[19] (
	.clk(clock),
	.d(\mepc[19]~17_combout ),
	.asdata(\_T_244[19]~31_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_19),
	.prn(vcc));
defparam \mepc[19] .is_wysiwyg = "true";
defparam \mepc[19] .power_up = "low";

dffeas \mepc[20] (
	.clk(clock),
	.d(\mepc[20]~18_combout ),
	.asdata(\_T_244[20]~33_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_20),
	.prn(vcc));
defparam \mepc[20] .is_wysiwyg = "true";
defparam \mepc[20] .power_up = "low";

dffeas \mepc[21] (
	.clk(clock),
	.d(\mepc[21]~19_combout ),
	.asdata(\_T_244[21]~35_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_21),
	.prn(vcc));
defparam \mepc[21] .is_wysiwyg = "true";
defparam \mepc[21] .power_up = "low";

dffeas \mepc[22] (
	.clk(clock),
	.d(\mepc[22]~20_combout ),
	.asdata(\_T_244[22]~37_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_22),
	.prn(vcc));
defparam \mepc[22] .is_wysiwyg = "true";
defparam \mepc[22] .power_up = "low";

dffeas \mepc[23] (
	.clk(clock),
	.d(\mepc[23]~21_combout ),
	.asdata(\_T_244[23]~39_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_23),
	.prn(vcc));
defparam \mepc[23] .is_wysiwyg = "true";
defparam \mepc[23] .power_up = "low";

dffeas \mepc[24] (
	.clk(clock),
	.d(\mepc[24]~22_combout ),
	.asdata(\_T_244[24]~41_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_24),
	.prn(vcc));
defparam \mepc[24] .is_wysiwyg = "true";
defparam \mepc[24] .power_up = "low";

dffeas \mepc[25] (
	.clk(clock),
	.d(\mepc[25]~23_combout ),
	.asdata(\_T_244[25]~43_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_25),
	.prn(vcc));
defparam \mepc[25] .is_wysiwyg = "true";
defparam \mepc[25] .power_up = "low";

dffeas \mepc[26] (
	.clk(clock),
	.d(\mepc[26]~24_combout ),
	.asdata(\_T_244[26]~45_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_26),
	.prn(vcc));
defparam \mepc[26] .is_wysiwyg = "true";
defparam \mepc[26] .power_up = "low";

dffeas \mepc[27] (
	.clk(clock),
	.d(\mepc[27]~25_combout ),
	.asdata(\_T_244[27]~47_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_27),
	.prn(vcc));
defparam \mepc[27] .is_wysiwyg = "true";
defparam \mepc[27] .power_up = "low";

dffeas \mepc[28] (
	.clk(clock),
	.d(\mepc[28]~26_combout ),
	.asdata(\_T_244[28]~49_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_28),
	.prn(vcc));
defparam \mepc[28] .is_wysiwyg = "true";
defparam \mepc[28] .power_up = "low";

dffeas \mepc[29] (
	.clk(clock),
	.d(\mepc[29]~27_combout ),
	.asdata(\_T_244[29]~51_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_29),
	.prn(vcc));
defparam \mepc[29] .is_wysiwyg = "true";
defparam \mepc[29] .power_up = "low";

dffeas \mepc[30] (
	.clk(clock),
	.d(\mepc[30]~28_combout ),
	.asdata(\_T_244[30]~53_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_30),
	.prn(vcc));
defparam \mepc[30] .is_wysiwyg = "true";
defparam \mepc[30] .power_up = "low";

dffeas \mepc[31] (
	.clk(clock),
	.d(\mepc[31]~29_combout ),
	.asdata(\_T_246[31]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(io_expt2),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_31),
	.prn(vcc));
defparam \mepc[31] .is_wysiwyg = "true";
defparam \mepc[31] .power_up = "low";

cyclone10lp_lcell_comb \io_expt~0 (
	.dataa(\mcause~4_combout ),
	.datab(\laddrInvalid~0_combout ),
	.datac(\saddrInvalid~0_combout ),
	.datad(\laddrInvalid~1_combout ),
	.cin(gnd),
	.combout(io_expt1),
	.cout());
defparam \io_expt~0 .lut_mask = 16'h08AA;
defparam \io_expt~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mcause[0]~6 (
	.dataa(\mcause[0]~5_combout ),
	.datab(read_latency_shift_reg_0),
	.datac(_T_3557),
	.datad(_T_3549),
	.cin(gnd),
	.combout(mcause_0),
	.cout());
defparam \mcause[0]~6 .lut_mask = 16'h0008;
defparam \mcause[0]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \isEcall~0 (
	.dataa(ex_csr_cmd_2),
	.datab(ex_csr_cmd_0),
	.datac(ex_csr_cmd_1),
	.datad(ex_csr_addr_8),
	.cin(gnd),
	.combout(isEcall),
	.cout());
defparam \isEcall~0 .lut_mask = 16'h0002;
defparam \isEcall~0 .sum_lutc_input = "datac";

dffeas \mepc[0] (
	.clk(clock),
	.d(\_GEN_204[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_0),
	.prn(vcc));
defparam \mepc[0] .is_wysiwyg = "true";
defparam \mepc[0] .power_up = "low";

cyclone10lp_lcell_comb io_expt(
	.dataa(io_expt1),
	.datab(gnd),
	.datac(gnd),
	.datad(isEcall),
	.cin(gnd),
	.combout(io_expt2),
	.cout());
defparam io_expt.lut_mask = 16'h00AA;
defparam io_expt.sum_lutc_input = "datac";

dffeas \mtvec[0] (
	.clk(clock),
	.d(\mtvec~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_0),
	.prn(vcc));
defparam \mtvec[0] .is_wysiwyg = "true";
defparam \mtvec[0] .power_up = "low";

dffeas \mepc[1] (
	.clk(clock),
	.d(\_GEN_204[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mepc[0]~30_combout ),
	.q(mepc_1),
	.prn(vcc));
defparam \mepc[1] .is_wysiwyg = "true";
defparam \mepc[1] .power_up = "low";

dffeas \mtvec[1] (
	.clk(clock),
	.d(\mtvec~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_1),
	.prn(vcc));
defparam \mtvec[1] .is_wysiwyg = "true";
defparam \mtvec[1] .power_up = "low";

cyclone10lp_lcell_comb \io_out[1]~16 (
	.dataa(\io_out[1]~7_combout ),
	.datab(\io_out[1]~9_combout ),
	.datac(\io_out[1]~11_combout ),
	.datad(\io_out[1]~15_combout ),
	.cin(gnd),
	.combout(io_out_1),
	.cout());
defparam \io_out[1]~16 .lut_mask = 16'hFFFE;
defparam \io_out[1]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[0]~24 (
	.dataa(\io_out[0]~21_combout ),
	.datab(\io_out[0]~23_combout ),
	.datac(\io_out[1]~14_combout ),
	.datad(\instreth[0]~q ),
	.cin(gnd),
	.combout(io_out_0),
	.cout());
defparam \io_out[0]~24 .lut_mask = 16'hFEEE;
defparam \io_out[0]~24 .sum_lutc_input = "datac";

dffeas \mtvec[2] (
	.clk(clock),
	.d(\mtvec~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_2),
	.prn(vcc));
defparam \mtvec[2] .is_wysiwyg = "true";
defparam \mtvec[2] .power_up = "low";

dffeas \mtvec[3] (
	.clk(clock),
	.d(\mtvec~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_3),
	.prn(vcc));
defparam \mtvec[3] .is_wysiwyg = "true";
defparam \mtvec[3] .power_up = "low";

dffeas \mtvec[4] (
	.clk(clock),
	.d(\mtvec~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_4),
	.prn(vcc));
defparam \mtvec[4] .is_wysiwyg = "true";
defparam \mtvec[4] .power_up = "low";

dffeas \mtvec[5] (
	.clk(clock),
	.d(\mtvec~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_5),
	.prn(vcc));
defparam \mtvec[5] .is_wysiwyg = "true";
defparam \mtvec[5] .power_up = "low";

dffeas \mtvec[6] (
	.clk(clock),
	.d(\mtvec~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_6),
	.prn(vcc));
defparam \mtvec[6] .is_wysiwyg = "true";
defparam \mtvec[6] .power_up = "low";

dffeas \mtvec[7] (
	.clk(clock),
	.d(\mtvec~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_7),
	.prn(vcc));
defparam \mtvec[7] .is_wysiwyg = "true";
defparam \mtvec[7] .power_up = "low";

dffeas \mtvec[8] (
	.clk(clock),
	.d(\mtvec~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_8),
	.prn(vcc));
defparam \mtvec[8] .is_wysiwyg = "true";
defparam \mtvec[8] .power_up = "low";

dffeas \mtvec[9] (
	.clk(clock),
	.d(\mtvec~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_9),
	.prn(vcc));
defparam \mtvec[9] .is_wysiwyg = "true";
defparam \mtvec[9] .power_up = "low";

dffeas \mtvec[10] (
	.clk(clock),
	.d(\mtvec~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_10),
	.prn(vcc));
defparam \mtvec[10] .is_wysiwyg = "true";
defparam \mtvec[10] .power_up = "low";

dffeas \mtvec[11] (
	.clk(clock),
	.d(\mtvec~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_11),
	.prn(vcc));
defparam \mtvec[11] .is_wysiwyg = "true";
defparam \mtvec[11] .power_up = "low";

dffeas \mtvec[12] (
	.clk(clock),
	.d(\mtvec~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_12),
	.prn(vcc));
defparam \mtvec[12] .is_wysiwyg = "true";
defparam \mtvec[12] .power_up = "low";

dffeas \mtvec[13] (
	.clk(clock),
	.d(\mtvec~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_13),
	.prn(vcc));
defparam \mtvec[13] .is_wysiwyg = "true";
defparam \mtvec[13] .power_up = "low";

dffeas \mtvec[14] (
	.clk(clock),
	.d(\mtvec~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_14),
	.prn(vcc));
defparam \mtvec[14] .is_wysiwyg = "true";
defparam \mtvec[14] .power_up = "low";

dffeas \mtvec[15] (
	.clk(clock),
	.d(\mtvec~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_15),
	.prn(vcc));
defparam \mtvec[15] .is_wysiwyg = "true";
defparam \mtvec[15] .power_up = "low";

dffeas \mtvec[16] (
	.clk(clock),
	.d(\mtvec~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_16),
	.prn(vcc));
defparam \mtvec[16] .is_wysiwyg = "true";
defparam \mtvec[16] .power_up = "low";

dffeas \mtvec[17] (
	.clk(clock),
	.d(\mtvec~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_17),
	.prn(vcc));
defparam \mtvec[17] .is_wysiwyg = "true";
defparam \mtvec[17] .power_up = "low";

dffeas \mtvec[18] (
	.clk(clock),
	.d(\mtvec~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_18),
	.prn(vcc));
defparam \mtvec[18] .is_wysiwyg = "true";
defparam \mtvec[18] .power_up = "low";

dffeas \mtvec[19] (
	.clk(clock),
	.d(\mtvec~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_19),
	.prn(vcc));
defparam \mtvec[19] .is_wysiwyg = "true";
defparam \mtvec[19] .power_up = "low";

dffeas \mtvec[20] (
	.clk(clock),
	.d(\mtvec~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_20),
	.prn(vcc));
defparam \mtvec[20] .is_wysiwyg = "true";
defparam \mtvec[20] .power_up = "low";

dffeas \mtvec[21] (
	.clk(clock),
	.d(\mtvec~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_21),
	.prn(vcc));
defparam \mtvec[21] .is_wysiwyg = "true";
defparam \mtvec[21] .power_up = "low";

dffeas \mtvec[22] (
	.clk(clock),
	.d(\mtvec~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_22),
	.prn(vcc));
defparam \mtvec[22] .is_wysiwyg = "true";
defparam \mtvec[22] .power_up = "low";

dffeas \mtvec[23] (
	.clk(clock),
	.d(\mtvec~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_23),
	.prn(vcc));
defparam \mtvec[23] .is_wysiwyg = "true";
defparam \mtvec[23] .power_up = "low";

dffeas \mtvec[24] (
	.clk(clock),
	.d(\mtvec~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_24),
	.prn(vcc));
defparam \mtvec[24] .is_wysiwyg = "true";
defparam \mtvec[24] .power_up = "low";

dffeas \mtvec[25] (
	.clk(clock),
	.d(\mtvec~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_25),
	.prn(vcc));
defparam \mtvec[25] .is_wysiwyg = "true";
defparam \mtvec[25] .power_up = "low";

dffeas \mtvec[26] (
	.clk(clock),
	.d(\mtvec~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_26),
	.prn(vcc));
defparam \mtvec[26] .is_wysiwyg = "true";
defparam \mtvec[26] .power_up = "low";

dffeas \mtvec[27] (
	.clk(clock),
	.d(\mtvec~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_27),
	.prn(vcc));
defparam \mtvec[27] .is_wysiwyg = "true";
defparam \mtvec[27] .power_up = "low";

dffeas \mtvec[28] (
	.clk(clock),
	.d(\mtvec~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_28),
	.prn(vcc));
defparam \mtvec[28] .is_wysiwyg = "true";
defparam \mtvec[28] .power_up = "low";

dffeas \mtvec[29] (
	.clk(clock),
	.d(\mtvec~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_29),
	.prn(vcc));
defparam \mtvec[29] .is_wysiwyg = "true";
defparam \mtvec[29] .power_up = "low";

dffeas \mtvec[30] (
	.clk(clock),
	.d(\mtvec~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_30),
	.prn(vcc));
defparam \mtvec[30] .is_wysiwyg = "true";
defparam \mtvec[30] .power_up = "low";

dffeas \mtvec[31] (
	.clk(clock),
	.d(\mtvec~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtvec[5]~1_combout ),
	.q(mtvec_31),
	.prn(vcc));
defparam \mtvec[31] .is_wysiwyg = "true";
defparam \mtvec[31] .power_up = "low";

cyclone10lp_lcell_comb \io_out[28]~31 (
	.dataa(\io_out[28]~29_combout ),
	.datab(\io_out[28]~30_combout ),
	.datac(\io_out[1]~12_combout ),
	.datad(\timeh[28]~q ),
	.cin(gnd),
	.combout(io_out_28),
	.cout());
defparam \io_out[28]~31 .lut_mask = 16'hFEEE;
defparam \io_out[28]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[29]~36 (
	.dataa(\io_out[29]~32_combout ),
	.datab(\io_out[29]~33_combout ),
	.datac(\io_out[29]~34_combout ),
	.datad(\io_out[29]~35_combout ),
	.cin(gnd),
	.combout(io_out_29),
	.cout());
defparam \io_out[29]~36 .lut_mask = 16'hFFFE;
defparam \io_out[29]~36 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[29]~37 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[29]~q ),
	.datad(\timeh[29]~q ),
	.cin(gnd),
	.combout(io_out_291),
	.cout());
defparam \io_out[29]~37 .lut_mask = 16'hEAC0;
defparam \io_out[29]~37 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[30]~45 (
	.dataa(\io_out[30]~41_combout ),
	.datab(\io_out[30]~42_combout ),
	.datac(\io_out[30]~43_combout ),
	.datad(\io_out[30]~44_combout ),
	.cin(gnd),
	.combout(io_out_30),
	.cout());
defparam \io_out[30]~45 .lut_mask = 16'hFFFE;
defparam \io_out[30]~45 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[31]~52 (
	.dataa(\io_out[31]~50_combout ),
	.datab(\io_out[31]~51_combout ),
	.datac(\io_out[1]~14_combout ),
	.datad(\instreth[31]~q ),
	.cin(gnd),
	.combout(io_out_31),
	.cout());
defparam \io_out[31]~52 .lut_mask = 16'hFEEE;
defparam \io_out[31]~52 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[8]~59 (
	.dataa(\io_out[8]~55_combout ),
	.datab(\io_out[8]~56_combout ),
	.datac(\io_out[8]~57_combout ),
	.datad(\io_out[8]~58_combout ),
	.cin(gnd),
	.combout(io_out_8),
	.cout());
defparam \io_out[8]~59 .lut_mask = 16'hFFFE;
defparam \io_out[8]~59 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[9]~66 (
	.dataa(\io_out[9]~60_combout ),
	.datab(\io_out[9]~61_combout ),
	.datac(\io_out[9]~64_combout ),
	.datad(\io_out[9]~65_combout ),
	.cin(gnd),
	.combout(io_out_9),
	.cout());
defparam \io_out[9]~66 .lut_mask = 16'hFFFE;
defparam \io_out[9]~66 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[10]~72 (
	.dataa(\io_out[10]~68_combout ),
	.datab(\io_out[10]~69_combout ),
	.datac(\io_out[10]~70_combout ),
	.datad(\io_out[10]~71_combout ),
	.cin(gnd),
	.combout(io_out_10),
	.cout());
defparam \io_out[10]~72 .lut_mask = 16'hFFFE;
defparam \io_out[10]~72 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[11]~79 (
	.dataa(\io_out[11]~73_combout ),
	.datab(\io_out[11]~74_combout ),
	.datac(\io_out[11]~77_combout ),
	.datad(\io_out[11]~78_combout ),
	.cin(gnd),
	.combout(io_out_11),
	.cout());
defparam \io_out[11]~79 .lut_mask = 16'hFFFE;
defparam \io_out[11]~79 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[12]~86 (
	.dataa(\io_out[12]~82_combout ),
	.datab(\io_out[12]~83_combout ),
	.datac(\io_out[12]~84_combout ),
	.datad(\io_out[12]~85_combout ),
	.cin(gnd),
	.combout(io_out_12),
	.cout());
defparam \io_out[12]~86 .lut_mask = 16'hFFFE;
defparam \io_out[12]~86 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[13]~93 (
	.dataa(\io_out[13]~91_combout ),
	.datab(\io_out[13]~92_combout ),
	.datac(\io_out[1]~12_combout ),
	.datad(\timeh[13]~q ),
	.cin(gnd),
	.combout(io_out_13),
	.cout());
defparam \io_out[13]~93 .lut_mask = 16'hFEEE;
defparam \io_out[13]~93 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[14]~100 (
	.dataa(\io_out[14]~96_combout ),
	.datab(\io_out[14]~97_combout ),
	.datac(\io_out[14]~98_combout ),
	.datad(\io_out[14]~99_combout ),
	.cin(gnd),
	.combout(io_out_14),
	.cout());
defparam \io_out[14]~100 .lut_mask = 16'hFFFE;
defparam \io_out[14]~100 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[15]~107 (
	.dataa(\io_out[15]~101_combout ),
	.datab(\io_out[15]~102_combout ),
	.datac(\io_out[15]~105_combout ),
	.datad(\io_out[15]~106_combout ),
	.cin(gnd),
	.combout(io_out_15),
	.cout());
defparam \io_out[15]~107 .lut_mask = 16'hFFFE;
defparam \io_out[15]~107 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[16]~114 (
	.dataa(\io_out[16]~110_combout ),
	.datab(\io_out[16]~111_combout ),
	.datac(\io_out[16]~112_combout ),
	.datad(\io_out[16]~113_combout ),
	.cin(gnd),
	.combout(io_out_16),
	.cout());
defparam \io_out[16]~114 .lut_mask = 16'hFFFE;
defparam \io_out[16]~114 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[17]~121 (
	.dataa(\io_out[17]~117_combout ),
	.datab(\io_out[17]~118_combout ),
	.datac(\io_out[17]~119_combout ),
	.datad(\io_out[17]~120_combout ),
	.cin(gnd),
	.combout(io_out_17),
	.cout());
defparam \io_out[17]~121 .lut_mask = 16'hFFFE;
defparam \io_out[17]~121 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[18]~128 (
	.dataa(\io_out[18]~126_combout ),
	.datab(\io_out[18]~127_combout ),
	.datac(\io_out[1]~12_combout ),
	.datad(\timeh[18]~q ),
	.cin(gnd),
	.combout(io_out_18),
	.cout());
defparam \io_out[18]~128 .lut_mask = 16'hFEEE;
defparam \io_out[18]~128 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[19]~135 (
	.dataa(\io_out[19]~129_combout ),
	.datab(\io_out[19]~130_combout ),
	.datac(\io_out[19]~133_combout ),
	.datad(\io_out[19]~134_combout ),
	.cin(gnd),
	.combout(io_out_19),
	.cout());
defparam \io_out[19]~135 .lut_mask = 16'hFFFE;
defparam \io_out[19]~135 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[4]~142 (
	.dataa(\io_out[4]~136_combout ),
	.datab(\io_out[4]~137_combout ),
	.datac(\io_out[4]~140_combout ),
	.datad(\io_out[4]~141_combout ),
	.cin(gnd),
	.combout(io_out_4),
	.cout());
defparam \io_out[4]~142 .lut_mask = 16'hFFFE;
defparam \io_out[4]~142 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[2]~150 (
	.dataa(\io_out[2]~145_combout ),
	.datab(\io_out[2]~146_combout ),
	.datac(\io_out[2]~147_combout ),
	.datad(\io_out[2]~149_combout ),
	.cin(gnd),
	.combout(io_out_2),
	.cout());
defparam \io_out[2]~150 .lut_mask = 16'hFFFE;
defparam \io_out[2]~150 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[3]~159 (
	.dataa(\io_out[3]~153_combout ),
	.datab(\io_out[3]~154_combout ),
	.datac(\io_out[3]~155_combout ),
	.datad(\io_out[3]~158_combout ),
	.cin(gnd),
	.combout(io_out_3),
	.cout());
defparam \io_out[3]~159 .lut_mask = 16'hFFFE;
defparam \io_out[3]~159 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[5]~166 (
	.dataa(\io_out[5]~160_combout ),
	.datab(\io_out[5]~161_combout ),
	.datac(\io_out[5]~164_combout ),
	.datad(\io_out[5]~165_combout ),
	.cin(gnd),
	.combout(io_out_5),
	.cout());
defparam \io_out[5]~166 .lut_mask = 16'hFFFE;
defparam \io_out[5]~166 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[6]~173 (
	.dataa(\io_out[6]~167_combout ),
	.datab(\io_out[6]~168_combout ),
	.datac(\io_out[6]~171_combout ),
	.datad(\io_out[6]~172_combout ),
	.cin(gnd),
	.combout(io_out_6),
	.cout());
defparam \io_out[6]~173 .lut_mask = 16'hFFFE;
defparam \io_out[6]~173 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[7]~181 (
	.dataa(\io_out[7]~179_combout ),
	.datab(\io_out[7]~180_combout ),
	.datac(\io_out[1]~14_combout ),
	.datad(\instreth[7]~q ),
	.cin(gnd),
	.combout(io_out_7),
	.cout());
defparam \io_out[7]~181 .lut_mask = 16'hFEEE;
defparam \io_out[7]~181 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[20]~188 (
	.dataa(\io_out[20]~184_combout ),
	.datab(\io_out[20]~185_combout ),
	.datac(\io_out[20]~186_combout ),
	.datad(\io_out[20]~187_combout ),
	.cin(gnd),
	.combout(io_out_20),
	.cout());
defparam \io_out[20]~188 .lut_mask = 16'hFFFE;
defparam \io_out[20]~188 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[21]~193 (
	.dataa(\io_out[21]~189_combout ),
	.datab(\io_out[21]~190_combout ),
	.datac(\io_out[21]~191_combout ),
	.datad(\io_out[21]~192_combout ),
	.cin(gnd),
	.combout(io_out_21),
	.cout());
defparam \io_out[21]~193 .lut_mask = 16'hFFFE;
defparam \io_out[21]~193 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[21]~194 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[21]~q ),
	.datad(\timeh[21]~q ),
	.cin(gnd),
	.combout(io_out_211),
	.cout());
defparam \io_out[21]~194 .lut_mask = 16'hEAC0;
defparam \io_out[21]~194 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[22]~202 (
	.dataa(\io_out[22]~196_combout ),
	.datab(\io_out[22]~197_combout ),
	.datac(\io_out[22]~200_combout ),
	.datad(\io_out[22]~201_combout ),
	.cin(gnd),
	.combout(io_out_22),
	.cout());
defparam \io_out[22]~202 .lut_mask = 16'hFFFE;
defparam \io_out[22]~202 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[23]~209 (
	.dataa(\io_out[23]~205_combout ),
	.datab(\io_out[23]~206_combout ),
	.datac(\io_out[23]~207_combout ),
	.datad(\io_out[23]~208_combout ),
	.cin(gnd),
	.combout(io_out_23),
	.cout());
defparam \io_out[23]~209 .lut_mask = 16'hFFFE;
defparam \io_out[23]~209 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[24]~216 (
	.dataa(\io_out[24]~210_combout ),
	.datab(\io_out[24]~211_combout ),
	.datac(\io_out[24]~214_combout ),
	.datad(\io_out[24]~215_combout ),
	.cin(gnd),
	.combout(io_out_24),
	.cout());
defparam \io_out[24]~216 .lut_mask = 16'hFFFE;
defparam \io_out[24]~216 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[25]~221 (
	.dataa(\io_out[25]~217_combout ),
	.datab(\io_out[25]~218_combout ),
	.datac(\io_out[25]~219_combout ),
	.datad(\io_out[25]~220_combout ),
	.cin(gnd),
	.combout(io_out_25),
	.cout());
defparam \io_out[25]~221 .lut_mask = 16'hFFFE;
defparam \io_out[25]~221 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[25]~222 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[25]~q ),
	.datad(\timeh[25]~q ),
	.cin(gnd),
	.combout(io_out_251),
	.cout());
defparam \io_out[25]~222 .lut_mask = 16'hEAC0;
defparam \io_out[25]~222 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[26]~230 (
	.dataa(\io_out[26]~226_combout ),
	.datab(\io_out[26]~227_combout ),
	.datac(\io_out[26]~228_combout ),
	.datad(\io_out[26]~229_combout ),
	.cin(gnd),
	.combout(io_out_26),
	.cout());
defparam \io_out[26]~230 .lut_mask = 16'hFFFE;
defparam \io_out[26]~230 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[27]~235 (
	.dataa(\io_out[27]~231_combout ),
	.datab(\io_out[27]~232_combout ),
	.datac(\io_out[27]~233_combout ),
	.datad(\io_out[27]~234_combout ),
	.cin(gnd),
	.combout(io_out_27),
	.cout());
defparam \io_out[27]~235 .lut_mask = 16'hFFFE;
defparam \io_out[27]~235 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[27]~236 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[27]~q ),
	.datad(\timeh[27]~q ),
	.cin(gnd),
	.combout(io_out_271),
	.cout());
defparam \io_out[27]~236 .lut_mask = 16'hEAC0;
defparam \io_out[27]~236 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~3 (
	.dataa(ex_pc_2),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~3_combout ),
	.cout());
defparam \pre_mepc~3 .lut_mask = 16'h8888;
defparam \pre_mepc~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc[28]~1 (
	.dataa(ex_j_check),
	.datab(ex_b_check),
	.datac(gnd),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\pre_mepc[28]~1_combout ),
	.cout());
defparam \pre_mepc[28]~1 .lut_mask = 16'hEEFF;
defparam \pre_mepc[28]~1 .sum_lutc_input = "datac";

dffeas \pre_mepc[2] (
	.clk(clock),
	.d(\pre_mepc~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[2]~q ),
	.prn(vcc));
defparam \pre_mepc[2] .is_wysiwyg = "true";
defparam \pre_mepc[2] .power_up = "low";

cyclone10lp_lcell_comb \mepc[2]~0 (
	.dataa(ex_pc_2),
	.datab(\pre_mepc[2]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[2]~0_combout ),
	.cout());
defparam \mepc[2]~0 .lut_mask = 16'hAACC;
defparam \mepc[2]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_246[0]~0 (
	.dataa(gnd),
	.datab(ex_csr_cmd_0),
	.datac(ex_csr_cmd_1),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_246[0]~0_combout ),
	.cout());
defparam \_T_246[0]~0 .lut_mask = 16'h003C;
defparam \_T_246[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_246[2]~5 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_2),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_246[2]~5_combout ),
	.cout());
defparam \_T_246[2]~5 .lut_mask = 16'h002A;
defparam \_T_246[2]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_246[2]~6 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_2),
	.datac(\_T_246[2]~5_combout ),
	.datad(csr_io_in_2),
	.cin(gnd),
	.combout(\_T_246[2]~6_combout ),
	.cout());
defparam \_T_246[2]~6 .lut_mask = 16'hEAC0;
defparam \_T_246[2]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal19~0 (
	.dataa(gnd),
	.datab(ex_csr_addr_4),
	.datac(ex_csr_addr_3),
	.datad(ex_csr_addr_5),
	.cin(gnd),
	.combout(\Equal19~0_combout ),
	.cout());
defparam \Equal19~0 .lut_mask = 16'h0003;
defparam \Equal19~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal25~2 (
	.dataa(\Equal19~0_combout ),
	.datab(ex_csr_addr_2),
	.datac(ex_csr_addr_10),
	.datad(ex_csr_addr_11),
	.cin(gnd),
	.combout(\Equal25~2_combout ),
	.cout());
defparam \Equal25~2 .lut_mask = 16'h0002;
defparam \Equal25~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal16~0 (
	.dataa(ex_csr_addr_8),
	.datab(ex_csr_addr_9),
	.datac(gnd),
	.datad(ex_csr_addr_7),
	.cin(gnd),
	.combout(\Equal16~0_combout ),
	.cout());
defparam \Equal16~0 .lut_mask = 16'h0088;
defparam \Equal16~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal4~0 (
	.dataa(ex_csr_addr_0),
	.datab(gnd),
	.datac(gnd),
	.datad(ex_csr_addr_1),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
defparam \Equal4~0 .lut_mask = 16'h00AA;
defparam \Equal4~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal26~0 (
	.dataa(ex_csr_addr_6),
	.datab(\Equal25~2_combout ),
	.datac(\Equal16~0_combout ),
	.datad(\Equal4~0_combout ),
	.cin(gnd),
	.combout(\Equal26~0_combout ),
	.cout());
defparam \Equal26~0 .lut_mask = 16'h8000;
defparam \Equal26~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb wen(
	.dataa(ex_csr_cmd_0),
	.datab(ex_csr_cmd_1),
	.datac(ex_csr_cmd_2),
	.datad(Equal59),
	.cin(gnd),
	.combout(\wen~combout ),
	.cout());
defparam wen.lut_mask = 16'h02CE;
defparam wen.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mepc[0]~30 (
	.dataa(io_expt2),
	.datab(\Equal26~0_combout ),
	.datac(\wen~combout ),
	.datad(mcause_0),
	.cin(gnd),
	.combout(\mepc[0]~30_combout ),
	.cout());
defparam \mepc[0]~30 .lut_mask = 16'hD500;
defparam \mepc[0]~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~4 (
	.dataa(ex_pc_3),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~4_combout ),
	.cout());
defparam \pre_mepc~4 .lut_mask = 16'h8888;
defparam \pre_mepc~4 .sum_lutc_input = "datac";

dffeas \pre_mepc[3] (
	.clk(clock),
	.d(\pre_mepc~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[3]~q ),
	.prn(vcc));
defparam \pre_mepc[3] .is_wysiwyg = "true";
defparam \pre_mepc[3] .power_up = "low";

cyclone10lp_lcell_comb \mepc[3]~1 (
	.dataa(ex_pc_3),
	.datab(\pre_mepc[3]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[3]~1_combout ),
	.cout());
defparam \mepc[3]~1 .lut_mask = 16'hAACC;
defparam \mepc[3]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_246[3]~7 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_3),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_246[3]~7_combout ),
	.cout());
defparam \_T_246[3]~7 .lut_mask = 16'h002A;
defparam \_T_246[3]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_246[3]~8 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_3),
	.datac(\_T_246[3]~7_combout ),
	.datad(csr_io_in_3),
	.cin(gnd),
	.combout(\_T_246[3]~8_combout ),
	.cout());
defparam \_T_246[3]~8 .lut_mask = 16'hEAC0;
defparam \_T_246[3]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~5 (
	.dataa(ex_pc_4),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~5_combout ),
	.cout());
defparam \pre_mepc~5 .lut_mask = 16'h8888;
defparam \pre_mepc~5 .sum_lutc_input = "datac";

dffeas \pre_mepc[4] (
	.clk(clock),
	.d(\pre_mepc~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[4]~q ),
	.prn(vcc));
defparam \pre_mepc[4] .is_wysiwyg = "true";
defparam \pre_mepc[4] .power_up = "low";

cyclone10lp_lcell_comb \mepc[4]~2 (
	.dataa(ex_pc_4),
	.datab(\pre_mepc[4]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[4]~2_combout ),
	.cout());
defparam \mepc[4]~2 .lut_mask = 16'hAACC;
defparam \mepc[4]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[4]~0 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_4),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[4]~0_combout ),
	.cout());
defparam \_T_244[4]~0 .lut_mask = 16'h002A;
defparam \_T_244[4]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[4]~1 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_4),
	.datac(\_T_244[4]~0_combout ),
	.datad(csr_io_in_4),
	.cin(gnd),
	.combout(\_T_244[4]~1_combout ),
	.cout());
defparam \_T_244[4]~1 .lut_mask = 16'hEAC0;
defparam \_T_244[4]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~6 (
	.dataa(ex_pc_5),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~6_combout ),
	.cout());
defparam \pre_mepc~6 .lut_mask = 16'h8888;
defparam \pre_mepc~6 .sum_lutc_input = "datac";

dffeas \pre_mepc[5] (
	.clk(clock),
	.d(\pre_mepc~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[5]~q ),
	.prn(vcc));
defparam \pre_mepc[5] .is_wysiwyg = "true";
defparam \pre_mepc[5] .power_up = "low";

cyclone10lp_lcell_comb \mepc[5]~3 (
	.dataa(ex_pc_5),
	.datab(\pre_mepc[5]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[5]~3_combout ),
	.cout());
defparam \mepc[5]~3 .lut_mask = 16'hAACC;
defparam \mepc[5]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[5]~2 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_5),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[5]~2_combout ),
	.cout());
defparam \_T_244[5]~2 .lut_mask = 16'h002A;
defparam \_T_244[5]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[5]~3 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_5),
	.datac(\_T_244[5]~2_combout ),
	.datad(csr_io_in_5),
	.cin(gnd),
	.combout(\_T_244[5]~3_combout ),
	.cout());
defparam \_T_244[5]~3 .lut_mask = 16'hEAC0;
defparam \_T_244[5]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~7 (
	.dataa(ex_pc_6),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~7_combout ),
	.cout());
defparam \pre_mepc~7 .lut_mask = 16'h8888;
defparam \pre_mepc~7 .sum_lutc_input = "datac";

dffeas \pre_mepc[6] (
	.clk(clock),
	.d(\pre_mepc~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[6]~q ),
	.prn(vcc));
defparam \pre_mepc[6] .is_wysiwyg = "true";
defparam \pre_mepc[6] .power_up = "low";

cyclone10lp_lcell_comb \mepc[6]~4 (
	.dataa(ex_pc_6),
	.datab(\pre_mepc[6]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[6]~4_combout ),
	.cout());
defparam \mepc[6]~4 .lut_mask = 16'hAACC;
defparam \mepc[6]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[6]~4 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_6),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[6]~4_combout ),
	.cout());
defparam \_T_244[6]~4 .lut_mask = 16'h002A;
defparam \_T_244[6]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[6]~5 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_6),
	.datac(\_T_244[6]~4_combout ),
	.datad(csr_io_in_6),
	.cin(gnd),
	.combout(\_T_244[6]~5_combout ),
	.cout());
defparam \_T_244[6]~5 .lut_mask = 16'hEAC0;
defparam \_T_244[6]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~8 (
	.dataa(ex_pc_7),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~8_combout ),
	.cout());
defparam \pre_mepc~8 .lut_mask = 16'h8888;
defparam \pre_mepc~8 .sum_lutc_input = "datac";

dffeas \pre_mepc[7] (
	.clk(clock),
	.d(\pre_mepc~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[7]~q ),
	.prn(vcc));
defparam \pre_mepc[7] .is_wysiwyg = "true";
defparam \pre_mepc[7] .power_up = "low";

cyclone10lp_lcell_comb \mepc[7]~5 (
	.dataa(ex_pc_7),
	.datab(\pre_mepc[7]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[7]~5_combout ),
	.cout());
defparam \mepc[7]~5 .lut_mask = 16'hAACC;
defparam \mepc[7]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[7]~6 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_7),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[7]~6_combout ),
	.cout());
defparam \_T_244[7]~6 .lut_mask = 16'h002A;
defparam \_T_244[7]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[7]~7 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_7),
	.datac(\_T_244[7]~6_combout ),
	.datad(csr_io_in_7),
	.cin(gnd),
	.combout(\_T_244[7]~7_combout ),
	.cout());
defparam \_T_244[7]~7 .lut_mask = 16'hEAC0;
defparam \_T_244[7]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~9 (
	.dataa(ex_pc_8),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~9_combout ),
	.cout());
defparam \pre_mepc~9 .lut_mask = 16'h8888;
defparam \pre_mepc~9 .sum_lutc_input = "datac";

dffeas \pre_mepc[8] (
	.clk(clock),
	.d(\pre_mepc~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[8]~q ),
	.prn(vcc));
defparam \pre_mepc[8] .is_wysiwyg = "true";
defparam \pre_mepc[8] .power_up = "low";

cyclone10lp_lcell_comb \mepc[8]~6 (
	.dataa(ex_pc_8),
	.datab(\pre_mepc[8]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[8]~6_combout ),
	.cout());
defparam \mepc[8]~6 .lut_mask = 16'hAACC;
defparam \mepc[8]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[8]~8 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_8),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[8]~8_combout ),
	.cout());
defparam \_T_244[8]~8 .lut_mask = 16'h002A;
defparam \_T_244[8]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[8]~9 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_8),
	.datac(\_T_244[8]~8_combout ),
	.datad(csr_io_in_8),
	.cin(gnd),
	.combout(\_T_244[8]~9_combout ),
	.cout());
defparam \_T_244[8]~9 .lut_mask = 16'hEAC0;
defparam \_T_244[8]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~10 (
	.dataa(ex_pc_9),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~10_combout ),
	.cout());
defparam \pre_mepc~10 .lut_mask = 16'h8888;
defparam \pre_mepc~10 .sum_lutc_input = "datac";

dffeas \pre_mepc[9] (
	.clk(clock),
	.d(\pre_mepc~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[9]~q ),
	.prn(vcc));
defparam \pre_mepc[9] .is_wysiwyg = "true";
defparam \pre_mepc[9] .power_up = "low";

cyclone10lp_lcell_comb \mepc[9]~7 (
	.dataa(ex_pc_9),
	.datab(\pre_mepc[9]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[9]~7_combout ),
	.cout());
defparam \mepc[9]~7 .lut_mask = 16'hAACC;
defparam \mepc[9]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[9]~10 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_9),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[9]~10_combout ),
	.cout());
defparam \_T_244[9]~10 .lut_mask = 16'h002A;
defparam \_T_244[9]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[9]~11 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_9),
	.datac(\_T_244[9]~10_combout ),
	.datad(csr_io_in_9),
	.cin(gnd),
	.combout(\_T_244[9]~11_combout ),
	.cout());
defparam \_T_244[9]~11 .lut_mask = 16'hEAC0;
defparam \_T_244[9]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~11 (
	.dataa(ex_pc_10),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~11_combout ),
	.cout());
defparam \pre_mepc~11 .lut_mask = 16'h8888;
defparam \pre_mepc~11 .sum_lutc_input = "datac";

dffeas \pre_mepc[10] (
	.clk(clock),
	.d(\pre_mepc~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[10]~q ),
	.prn(vcc));
defparam \pre_mepc[10] .is_wysiwyg = "true";
defparam \pre_mepc[10] .power_up = "low";

cyclone10lp_lcell_comb \mepc[10]~8 (
	.dataa(ex_pc_10),
	.datab(\pre_mepc[10]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[10]~8_combout ),
	.cout());
defparam \mepc[10]~8 .lut_mask = 16'hAACC;
defparam \mepc[10]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[10]~12 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_10),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[10]~12_combout ),
	.cout());
defparam \_T_244[10]~12 .lut_mask = 16'h002A;
defparam \_T_244[10]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[10]~13 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_10),
	.datac(\_T_244[10]~12_combout ),
	.datad(csr_io_in_10),
	.cin(gnd),
	.combout(\_T_244[10]~13_combout ),
	.cout());
defparam \_T_244[10]~13 .lut_mask = 16'hEAC0;
defparam \_T_244[10]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~12 (
	.dataa(ex_pc_11),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~12_combout ),
	.cout());
defparam \pre_mepc~12 .lut_mask = 16'h8888;
defparam \pre_mepc~12 .sum_lutc_input = "datac";

dffeas \pre_mepc[11] (
	.clk(clock),
	.d(\pre_mepc~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[11]~q ),
	.prn(vcc));
defparam \pre_mepc[11] .is_wysiwyg = "true";
defparam \pre_mepc[11] .power_up = "low";

cyclone10lp_lcell_comb \mepc[11]~9 (
	.dataa(ex_pc_11),
	.datab(\pre_mepc[11]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[11]~9_combout ),
	.cout());
defparam \mepc[11]~9 .lut_mask = 16'hAACC;
defparam \mepc[11]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[11]~14 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_11),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[11]~14_combout ),
	.cout());
defparam \_T_244[11]~14 .lut_mask = 16'h002A;
defparam \_T_244[11]~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[11]~15 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_11),
	.datac(\_T_244[11]~14_combout ),
	.datad(csr_io_in_11),
	.cin(gnd),
	.combout(\_T_244[11]~15_combout ),
	.cout());
defparam \_T_244[11]~15 .lut_mask = 16'hEAC0;
defparam \_T_244[11]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~13 (
	.dataa(ex_pc_12),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~13_combout ),
	.cout());
defparam \pre_mepc~13 .lut_mask = 16'h8888;
defparam \pre_mepc~13 .sum_lutc_input = "datac";

dffeas \pre_mepc[12] (
	.clk(clock),
	.d(\pre_mepc~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[12]~q ),
	.prn(vcc));
defparam \pre_mepc[12] .is_wysiwyg = "true";
defparam \pre_mepc[12] .power_up = "low";

cyclone10lp_lcell_comb \mepc[12]~10 (
	.dataa(ex_pc_12),
	.datab(\pre_mepc[12]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[12]~10_combout ),
	.cout());
defparam \mepc[12]~10 .lut_mask = 16'hAACC;
defparam \mepc[12]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[12]~16 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_12),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[12]~16_combout ),
	.cout());
defparam \_T_244[12]~16 .lut_mask = 16'h002A;
defparam \_T_244[12]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[12]~17 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_12),
	.datac(\_T_244[12]~16_combout ),
	.datad(csr_io_in_12),
	.cin(gnd),
	.combout(\_T_244[12]~17_combout ),
	.cout());
defparam \_T_244[12]~17 .lut_mask = 16'hEAC0;
defparam \_T_244[12]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~14 (
	.dataa(ex_pc_13),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~14_combout ),
	.cout());
defparam \pre_mepc~14 .lut_mask = 16'h8888;
defparam \pre_mepc~14 .sum_lutc_input = "datac";

dffeas \pre_mepc[13] (
	.clk(clock),
	.d(\pre_mepc~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[13]~q ),
	.prn(vcc));
defparam \pre_mepc[13] .is_wysiwyg = "true";
defparam \pre_mepc[13] .power_up = "low";

cyclone10lp_lcell_comb \mepc[13]~11 (
	.dataa(ex_pc_13),
	.datab(\pre_mepc[13]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[13]~11_combout ),
	.cout());
defparam \mepc[13]~11 .lut_mask = 16'hAACC;
defparam \mepc[13]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[13]~18 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_13),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[13]~18_combout ),
	.cout());
defparam \_T_244[13]~18 .lut_mask = 16'h002A;
defparam \_T_244[13]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[13]~19 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_13),
	.datac(\_T_244[13]~18_combout ),
	.datad(csr_io_in_13),
	.cin(gnd),
	.combout(\_T_244[13]~19_combout ),
	.cout());
defparam \_T_244[13]~19 .lut_mask = 16'hEAC0;
defparam \_T_244[13]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~15 (
	.dataa(ex_pc_14),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~15_combout ),
	.cout());
defparam \pre_mepc~15 .lut_mask = 16'h8888;
defparam \pre_mepc~15 .sum_lutc_input = "datac";

dffeas \pre_mepc[14] (
	.clk(clock),
	.d(\pre_mepc~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[14]~q ),
	.prn(vcc));
defparam \pre_mepc[14] .is_wysiwyg = "true";
defparam \pre_mepc[14] .power_up = "low";

cyclone10lp_lcell_comb \mepc[14]~12 (
	.dataa(ex_pc_14),
	.datab(\pre_mepc[14]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[14]~12_combout ),
	.cout());
defparam \mepc[14]~12 .lut_mask = 16'hAACC;
defparam \mepc[14]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[14]~20 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_14),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[14]~20_combout ),
	.cout());
defparam \_T_244[14]~20 .lut_mask = 16'h002A;
defparam \_T_244[14]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[14]~21 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_14),
	.datac(\_T_244[14]~20_combout ),
	.datad(csr_io_in_14),
	.cin(gnd),
	.combout(\_T_244[14]~21_combout ),
	.cout());
defparam \_T_244[14]~21 .lut_mask = 16'hEAC0;
defparam \_T_244[14]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~16 (
	.dataa(ex_pc_15),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~16_combout ),
	.cout());
defparam \pre_mepc~16 .lut_mask = 16'h8888;
defparam \pre_mepc~16 .sum_lutc_input = "datac";

dffeas \pre_mepc[15] (
	.clk(clock),
	.d(\pre_mepc~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[15]~q ),
	.prn(vcc));
defparam \pre_mepc[15] .is_wysiwyg = "true";
defparam \pre_mepc[15] .power_up = "low";

cyclone10lp_lcell_comb \mepc[15]~13 (
	.dataa(ex_pc_15),
	.datab(\pre_mepc[15]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[15]~13_combout ),
	.cout());
defparam \mepc[15]~13 .lut_mask = 16'hAACC;
defparam \mepc[15]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[15]~22 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_15),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[15]~22_combout ),
	.cout());
defparam \_T_244[15]~22 .lut_mask = 16'h002A;
defparam \_T_244[15]~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[15]~23 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_15),
	.datac(\_T_244[15]~22_combout ),
	.datad(csr_io_in_15),
	.cin(gnd),
	.combout(\_T_244[15]~23_combout ),
	.cout());
defparam \_T_244[15]~23 .lut_mask = 16'hEAC0;
defparam \_T_244[15]~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~17 (
	.dataa(ex_pc_16),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~17_combout ),
	.cout());
defparam \pre_mepc~17 .lut_mask = 16'h8888;
defparam \pre_mepc~17 .sum_lutc_input = "datac";

dffeas \pre_mepc[16] (
	.clk(clock),
	.d(\pre_mepc~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[16]~q ),
	.prn(vcc));
defparam \pre_mepc[16] .is_wysiwyg = "true";
defparam \pre_mepc[16] .power_up = "low";

cyclone10lp_lcell_comb \mepc[16]~14 (
	.dataa(ex_pc_16),
	.datab(\pre_mepc[16]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[16]~14_combout ),
	.cout());
defparam \mepc[16]~14 .lut_mask = 16'hAACC;
defparam \mepc[16]~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[16]~24 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_16),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[16]~24_combout ),
	.cout());
defparam \_T_244[16]~24 .lut_mask = 16'h002A;
defparam \_T_244[16]~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[16]~25 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_16),
	.datac(\_T_244[16]~24_combout ),
	.datad(csr_io_in_16),
	.cin(gnd),
	.combout(\_T_244[16]~25_combout ),
	.cout());
defparam \_T_244[16]~25 .lut_mask = 16'hEAC0;
defparam \_T_244[16]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~18 (
	.dataa(ex_pc_17),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~18_combout ),
	.cout());
defparam \pre_mepc~18 .lut_mask = 16'h8888;
defparam \pre_mepc~18 .sum_lutc_input = "datac";

dffeas \pre_mepc[17] (
	.clk(clock),
	.d(\pre_mepc~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[17]~q ),
	.prn(vcc));
defparam \pre_mepc[17] .is_wysiwyg = "true";
defparam \pre_mepc[17] .power_up = "low";

cyclone10lp_lcell_comb \mepc[17]~15 (
	.dataa(ex_pc_17),
	.datab(\pre_mepc[17]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[17]~15_combout ),
	.cout());
defparam \mepc[17]~15 .lut_mask = 16'hAACC;
defparam \mepc[17]~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[17]~26 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_17),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[17]~26_combout ),
	.cout());
defparam \_T_244[17]~26 .lut_mask = 16'h002A;
defparam \_T_244[17]~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[17]~27 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_17),
	.datac(\_T_244[17]~26_combout ),
	.datad(csr_io_in_17),
	.cin(gnd),
	.combout(\_T_244[17]~27_combout ),
	.cout());
defparam \_T_244[17]~27 .lut_mask = 16'hEAC0;
defparam \_T_244[17]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~19 (
	.dataa(ex_pc_18),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~19_combout ),
	.cout());
defparam \pre_mepc~19 .lut_mask = 16'h8888;
defparam \pre_mepc~19 .sum_lutc_input = "datac";

dffeas \pre_mepc[18] (
	.clk(clock),
	.d(\pre_mepc~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[18]~q ),
	.prn(vcc));
defparam \pre_mepc[18] .is_wysiwyg = "true";
defparam \pre_mepc[18] .power_up = "low";

cyclone10lp_lcell_comb \mepc[18]~16 (
	.dataa(ex_pc_18),
	.datab(\pre_mepc[18]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[18]~16_combout ),
	.cout());
defparam \mepc[18]~16 .lut_mask = 16'hAACC;
defparam \mepc[18]~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[18]~28 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_18),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[18]~28_combout ),
	.cout());
defparam \_T_244[18]~28 .lut_mask = 16'h002A;
defparam \_T_244[18]~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[18]~29 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_18),
	.datac(\_T_244[18]~28_combout ),
	.datad(csr_io_in_18),
	.cin(gnd),
	.combout(\_T_244[18]~29_combout ),
	.cout());
defparam \_T_244[18]~29 .lut_mask = 16'hEAC0;
defparam \_T_244[18]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~20 (
	.dataa(ex_pc_19),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~20_combout ),
	.cout());
defparam \pre_mepc~20 .lut_mask = 16'h8888;
defparam \pre_mepc~20 .sum_lutc_input = "datac";

dffeas \pre_mepc[19] (
	.clk(clock),
	.d(\pre_mepc~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[19]~q ),
	.prn(vcc));
defparam \pre_mepc[19] .is_wysiwyg = "true";
defparam \pre_mepc[19] .power_up = "low";

cyclone10lp_lcell_comb \mepc[19]~17 (
	.dataa(ex_pc_19),
	.datab(\pre_mepc[19]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[19]~17_combout ),
	.cout());
defparam \mepc[19]~17 .lut_mask = 16'hAACC;
defparam \mepc[19]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[19]~30 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_19),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[19]~30_combout ),
	.cout());
defparam \_T_244[19]~30 .lut_mask = 16'h002A;
defparam \_T_244[19]~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[19]~31 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_19),
	.datac(\_T_244[19]~30_combout ),
	.datad(csr_io_in_19),
	.cin(gnd),
	.combout(\_T_244[19]~31_combout ),
	.cout());
defparam \_T_244[19]~31 .lut_mask = 16'hEAC0;
defparam \_T_244[19]~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~21 (
	.dataa(ex_pc_20),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~21_combout ),
	.cout());
defparam \pre_mepc~21 .lut_mask = 16'h8888;
defparam \pre_mepc~21 .sum_lutc_input = "datac";

dffeas \pre_mepc[20] (
	.clk(clock),
	.d(\pre_mepc~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[20]~q ),
	.prn(vcc));
defparam \pre_mepc[20] .is_wysiwyg = "true";
defparam \pre_mepc[20] .power_up = "low";

cyclone10lp_lcell_comb \mepc[20]~18 (
	.dataa(ex_pc_20),
	.datab(\pre_mepc[20]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[20]~18_combout ),
	.cout());
defparam \mepc[20]~18 .lut_mask = 16'hAACC;
defparam \mepc[20]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[20]~32 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_20),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[20]~32_combout ),
	.cout());
defparam \_T_244[20]~32 .lut_mask = 16'h002A;
defparam \_T_244[20]~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[20]~33 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_20),
	.datac(\_T_244[20]~32_combout ),
	.datad(csr_io_in_20),
	.cin(gnd),
	.combout(\_T_244[20]~33_combout ),
	.cout());
defparam \_T_244[20]~33 .lut_mask = 16'hEAC0;
defparam \_T_244[20]~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~22 (
	.dataa(ex_pc_21),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~22_combout ),
	.cout());
defparam \pre_mepc~22 .lut_mask = 16'h8888;
defparam \pre_mepc~22 .sum_lutc_input = "datac";

dffeas \pre_mepc[21] (
	.clk(clock),
	.d(\pre_mepc~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[21]~q ),
	.prn(vcc));
defparam \pre_mepc[21] .is_wysiwyg = "true";
defparam \pre_mepc[21] .power_up = "low";

cyclone10lp_lcell_comb \mepc[21]~19 (
	.dataa(ex_pc_21),
	.datab(\pre_mepc[21]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[21]~19_combout ),
	.cout());
defparam \mepc[21]~19 .lut_mask = 16'hAACC;
defparam \mepc[21]~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[21]~195 (
	.dataa(io_out_21),
	.datab(io_out_211),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[21]~195_combout ),
	.cout());
defparam \io_out[21]~195 .lut_mask = 16'hEEEE;
defparam \io_out[21]~195 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[21]~34 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_21),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[21]~34_combout ),
	.cout());
defparam \_T_244[21]~34 .lut_mask = 16'h002A;
defparam \_T_244[21]~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[21]~35 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(\io_out[21]~195_combout ),
	.datac(\_T_244[21]~34_combout ),
	.datad(csr_io_in_21),
	.cin(gnd),
	.combout(\_T_244[21]~35_combout ),
	.cout());
defparam \_T_244[21]~35 .lut_mask = 16'hEAC0;
defparam \_T_244[21]~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~23 (
	.dataa(ex_pc_22),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~23_combout ),
	.cout());
defparam \pre_mepc~23 .lut_mask = 16'h8888;
defparam \pre_mepc~23 .sum_lutc_input = "datac";

dffeas \pre_mepc[22] (
	.clk(clock),
	.d(\pre_mepc~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[22]~q ),
	.prn(vcc));
defparam \pre_mepc[22] .is_wysiwyg = "true";
defparam \pre_mepc[22] .power_up = "low";

cyclone10lp_lcell_comb \mepc[22]~20 (
	.dataa(ex_pc_22),
	.datab(\pre_mepc[22]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[22]~20_combout ),
	.cout());
defparam \mepc[22]~20 .lut_mask = 16'hAACC;
defparam \mepc[22]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[22]~36 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_22),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[22]~36_combout ),
	.cout());
defparam \_T_244[22]~36 .lut_mask = 16'h002A;
defparam \_T_244[22]~36 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[22]~37 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_22),
	.datac(\_T_244[22]~36_combout ),
	.datad(csr_io_in_22),
	.cin(gnd),
	.combout(\_T_244[22]~37_combout ),
	.cout());
defparam \_T_244[22]~37 .lut_mask = 16'hEAC0;
defparam \_T_244[22]~37 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~24 (
	.dataa(ex_pc_23),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~24_combout ),
	.cout());
defparam \pre_mepc~24 .lut_mask = 16'h8888;
defparam \pre_mepc~24 .sum_lutc_input = "datac";

dffeas \pre_mepc[23] (
	.clk(clock),
	.d(\pre_mepc~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[23]~q ),
	.prn(vcc));
defparam \pre_mepc[23] .is_wysiwyg = "true";
defparam \pre_mepc[23] .power_up = "low";

cyclone10lp_lcell_comb \mepc[23]~21 (
	.dataa(ex_pc_23),
	.datab(\pre_mepc[23]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[23]~21_combout ),
	.cout());
defparam \mepc[23]~21 .lut_mask = 16'hAACC;
defparam \mepc[23]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[23]~38 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_23),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[23]~38_combout ),
	.cout());
defparam \_T_244[23]~38 .lut_mask = 16'h002A;
defparam \_T_244[23]~38 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[23]~39 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_23),
	.datac(\_T_244[23]~38_combout ),
	.datad(csr_io_in_23),
	.cin(gnd),
	.combout(\_T_244[23]~39_combout ),
	.cout());
defparam \_T_244[23]~39 .lut_mask = 16'hEAC0;
defparam \_T_244[23]~39 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~25 (
	.dataa(ex_pc_24),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~25_combout ),
	.cout());
defparam \pre_mepc~25 .lut_mask = 16'h8888;
defparam \pre_mepc~25 .sum_lutc_input = "datac";

dffeas \pre_mepc[24] (
	.clk(clock),
	.d(\pre_mepc~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[24]~q ),
	.prn(vcc));
defparam \pre_mepc[24] .is_wysiwyg = "true";
defparam \pre_mepc[24] .power_up = "low";

cyclone10lp_lcell_comb \mepc[24]~22 (
	.dataa(ex_pc_24),
	.datab(\pre_mepc[24]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[24]~22_combout ),
	.cout());
defparam \mepc[24]~22 .lut_mask = 16'hAACC;
defparam \mepc[24]~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[24]~40 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_24),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[24]~40_combout ),
	.cout());
defparam \_T_244[24]~40 .lut_mask = 16'h002A;
defparam \_T_244[24]~40 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[24]~41 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_24),
	.datac(\_T_244[24]~40_combout ),
	.datad(csr_io_in_24),
	.cin(gnd),
	.combout(\_T_244[24]~41_combout ),
	.cout());
defparam \_T_244[24]~41 .lut_mask = 16'hEAC0;
defparam \_T_244[24]~41 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~26 (
	.dataa(ex_pc_25),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~26_combout ),
	.cout());
defparam \pre_mepc~26 .lut_mask = 16'h8888;
defparam \pre_mepc~26 .sum_lutc_input = "datac";

dffeas \pre_mepc[25] (
	.clk(clock),
	.d(\pre_mepc~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[25]~q ),
	.prn(vcc));
defparam \pre_mepc[25] .is_wysiwyg = "true";
defparam \pre_mepc[25] .power_up = "low";

cyclone10lp_lcell_comb \mepc[25]~23 (
	.dataa(ex_pc_25),
	.datab(\pre_mepc[25]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[25]~23_combout ),
	.cout());
defparam \mepc[25]~23 .lut_mask = 16'hAACC;
defparam \mepc[25]~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[25]~223 (
	.dataa(io_out_25),
	.datab(io_out_251),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[25]~223_combout ),
	.cout());
defparam \io_out[25]~223 .lut_mask = 16'hEEEE;
defparam \io_out[25]~223 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[25]~42 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_25),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[25]~42_combout ),
	.cout());
defparam \_T_244[25]~42 .lut_mask = 16'h002A;
defparam \_T_244[25]~42 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[25]~43 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(\io_out[25]~223_combout ),
	.datac(\_T_244[25]~42_combout ),
	.datad(csr_io_in_25),
	.cin(gnd),
	.combout(\_T_244[25]~43_combout ),
	.cout());
defparam \_T_244[25]~43 .lut_mask = 16'hEAC0;
defparam \_T_244[25]~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~27 (
	.dataa(ex_pc_26),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~27_combout ),
	.cout());
defparam \pre_mepc~27 .lut_mask = 16'h8888;
defparam \pre_mepc~27 .sum_lutc_input = "datac";

dffeas \pre_mepc[26] (
	.clk(clock),
	.d(\pre_mepc~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[26]~q ),
	.prn(vcc));
defparam \pre_mepc[26] .is_wysiwyg = "true";
defparam \pre_mepc[26] .power_up = "low";

cyclone10lp_lcell_comb \mepc[26]~24 (
	.dataa(ex_pc_26),
	.datab(\pre_mepc[26]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[26]~24_combout ),
	.cout());
defparam \mepc[26]~24 .lut_mask = 16'hAACC;
defparam \mepc[26]~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[26]~44 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_26),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[26]~44_combout ),
	.cout());
defparam \_T_244[26]~44 .lut_mask = 16'h002A;
defparam \_T_244[26]~44 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[26]~45 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_26),
	.datac(\_T_244[26]~44_combout ),
	.datad(csr_io_in_26),
	.cin(gnd),
	.combout(\_T_244[26]~45_combout ),
	.cout());
defparam \_T_244[26]~45 .lut_mask = 16'hEAC0;
defparam \_T_244[26]~45 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~28 (
	.dataa(ex_pc_27),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~28_combout ),
	.cout());
defparam \pre_mepc~28 .lut_mask = 16'h8888;
defparam \pre_mepc~28 .sum_lutc_input = "datac";

dffeas \pre_mepc[27] (
	.clk(clock),
	.d(\pre_mepc~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[27]~q ),
	.prn(vcc));
defparam \pre_mepc[27] .is_wysiwyg = "true";
defparam \pre_mepc[27] .power_up = "low";

cyclone10lp_lcell_comb \mepc[27]~25 (
	.dataa(ex_pc_27),
	.datab(\pre_mepc[27]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[27]~25_combout ),
	.cout());
defparam \mepc[27]~25 .lut_mask = 16'hAACC;
defparam \mepc[27]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[27]~237 (
	.dataa(io_out_27),
	.datab(io_out_271),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[27]~237_combout ),
	.cout());
defparam \io_out[27]~237 .lut_mask = 16'hEEEE;
defparam \io_out[27]~237 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[27]~46 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_27),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[27]~46_combout ),
	.cout());
defparam \_T_244[27]~46 .lut_mask = 16'h002A;
defparam \_T_244[27]~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[27]~47 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(\io_out[27]~237_combout ),
	.datac(\_T_244[27]~46_combout ),
	.datad(csr_io_in_27),
	.cin(gnd),
	.combout(\_T_244[27]~47_combout ),
	.cout());
defparam \_T_244[27]~47 .lut_mask = 16'hEAC0;
defparam \_T_244[27]~47 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~29 (
	.dataa(ex_pc_28),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~29_combout ),
	.cout());
defparam \pre_mepc~29 .lut_mask = 16'h8888;
defparam \pre_mepc~29 .sum_lutc_input = "datac";

dffeas \pre_mepc[28] (
	.clk(clock),
	.d(\pre_mepc~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[28]~q ),
	.prn(vcc));
defparam \pre_mepc[28] .is_wysiwyg = "true";
defparam \pre_mepc[28] .power_up = "low";

cyclone10lp_lcell_comb \mepc[28]~26 (
	.dataa(ex_pc_28),
	.datab(\pre_mepc[28]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[28]~26_combout ),
	.cout());
defparam \mepc[28]~26 .lut_mask = 16'hAACC;
defparam \mepc[28]~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[28]~48 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_28),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[28]~48_combout ),
	.cout());
defparam \_T_244[28]~48 .lut_mask = 16'h002A;
defparam \_T_244[28]~48 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[28]~49 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_28),
	.datac(\_T_244[28]~48_combout ),
	.datad(csr_io_in_28),
	.cin(gnd),
	.combout(\_T_244[28]~49_combout ),
	.cout());
defparam \_T_244[28]~49 .lut_mask = 16'hEAC0;
defparam \_T_244[28]~49 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~30 (
	.dataa(ex_pc_29),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~30_combout ),
	.cout());
defparam \pre_mepc~30 .lut_mask = 16'h8888;
defparam \pre_mepc~30 .sum_lutc_input = "datac";

dffeas \pre_mepc[29] (
	.clk(clock),
	.d(\pre_mepc~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[29]~q ),
	.prn(vcc));
defparam \pre_mepc[29] .is_wysiwyg = "true";
defparam \pre_mepc[29] .power_up = "low";

cyclone10lp_lcell_comb \mepc[29]~27 (
	.dataa(ex_pc_29),
	.datab(\pre_mepc[29]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[29]~27_combout ),
	.cout());
defparam \mepc[29]~27 .lut_mask = 16'hAACC;
defparam \mepc[29]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[29]~38 (
	.dataa(io_out_29),
	.datab(io_out_291),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[29]~38_combout ),
	.cout());
defparam \io_out[29]~38 .lut_mask = 16'hEEEE;
defparam \io_out[29]~38 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[29]~50 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_29),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[29]~50_combout ),
	.cout());
defparam \_T_244[29]~50 .lut_mask = 16'h002A;
defparam \_T_244[29]~50 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[29]~51 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(\io_out[29]~38_combout ),
	.datac(\_T_244[29]~50_combout ),
	.datad(csr_io_in_29),
	.cin(gnd),
	.combout(\_T_244[29]~51_combout ),
	.cout());
defparam \_T_244[29]~51 .lut_mask = 16'hEAC0;
defparam \_T_244[29]~51 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~31 (
	.dataa(ex_pc_30),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~31_combout ),
	.cout());
defparam \pre_mepc~31 .lut_mask = 16'h8888;
defparam \pre_mepc~31 .sum_lutc_input = "datac";

dffeas \pre_mepc[30] (
	.clk(clock),
	.d(\pre_mepc~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[30]~q ),
	.prn(vcc));
defparam \pre_mepc[30] .is_wysiwyg = "true";
defparam \pre_mepc[30] .power_up = "low";

cyclone10lp_lcell_comb \mepc[30]~28 (
	.dataa(ex_pc_30),
	.datab(\pre_mepc[30]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[30]~28_combout ),
	.cout());
defparam \mepc[30]~28 .lut_mask = 16'hAACC;
defparam \mepc[30]~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[30]~52 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_30),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_244[30]~52_combout ),
	.cout());
defparam \_T_244[30]~52 .lut_mask = 16'h002A;
defparam \_T_244[30]~52 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_244[30]~53 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_30),
	.datac(\_T_244[30]~52_combout ),
	.datad(csr_io_in_30),
	.cin(gnd),
	.combout(\_T_244[30]~53_combout ),
	.cout());
defparam \_T_244[30]~53 .lut_mask = 16'hEAC0;
defparam \_T_244[30]~53 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~32 (
	.dataa(ex_pc_31),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~32_combout ),
	.cout());
defparam \pre_mepc~32 .lut_mask = 16'h8888;
defparam \pre_mepc~32 .sum_lutc_input = "datac";

dffeas \pre_mepc[31] (
	.clk(clock),
	.d(\pre_mepc~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[31]~q ),
	.prn(vcc));
defparam \pre_mepc[31] .is_wysiwyg = "true";
defparam \pre_mepc[31] .power_up = "low";

cyclone10lp_lcell_comb \mepc[31]~29 (
	.dataa(ex_pc_31),
	.datab(\pre_mepc[31]~q ),
	.datac(gnd),
	.datad(Equal56),
	.cin(gnd),
	.combout(\mepc[31]~29_combout ),
	.cout());
defparam \mepc[31]~29 .lut_mask = 16'hAACC;
defparam \mepc[31]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_246[31]~9 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_31),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_246[31]~9_combout ),
	.cout());
defparam \_T_246[31]~9 .lut_mask = 16'h002A;
defparam \_T_246[31]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_246[31]~10 (
	.dataa(\_T_246[0]~0_combout ),
	.datab(io_out_31),
	.datac(\_T_246[31]~9_combout ),
	.datad(csr_io_in_31),
	.cin(gnd),
	.combout(\_T_246[31]~10_combout ),
	.cout());
defparam \_T_246[31]~10 .lut_mask = 16'hEAC0;
defparam \_T_246[31]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \isIllegal~0 (
	.dataa(Equal561),
	.datab(ex_ctrl_legal),
	.datac(gnd),
	.datad(inst_kill),
	.cin(gnd),
	.combout(\isIllegal~0_combout ),
	.cout());
defparam \isIllegal~0 .lut_mask = 16'hEEFF;
defparam \isIllegal~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \iaddrInvalid_j~0 (
	.dataa(csr_io_alu_op1_1),
	.datab(csr_io_alu_op2_1),
	.datac(csr_io_alu_op2_0),
	.datad(csr_io_alu_op1_0),
	.cin(gnd),
	.combout(\iaddrInvalid_j~0_combout ),
	.cout());
defparam \iaddrInvalid_j~0 .lut_mask = 16'h9FF6;
defparam \iaddrInvalid_j~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mcause~4 (
	.dataa(Equal56),
	.datab(\isIllegal~0_combout ),
	.datac(ex_j_check),
	.datad(\iaddrInvalid_j~0_combout ),
	.cin(gnd),
	.combout(\mcause~4_combout ),
	.cout());
defparam \mcause~4 .lut_mask = 16'h0888;
defparam \mcause~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \laddrInvalid~0 (
	.dataa(ex_ctrl_mask_type_0),
	.datab(ex_ctrl_mask_type_2),
	.datac(gnd),
	.datad(ex_ctrl_mem_wr01),
	.cin(gnd),
	.combout(\laddrInvalid~0_combout ),
	.cout());
defparam \laddrInvalid~0 .lut_mask = 16'h88FF;
defparam \laddrInvalid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \saddrInvalid~0 (
	.dataa(ex_ctrl_imm_type001),
	.datab(gnd),
	.datac(gnd),
	.datad(ex_ctrl_mask_type_2),
	.cin(gnd),
	.combout(\saddrInvalid~0_combout ),
	.cout());
defparam \saddrInvalid~0 .lut_mask = 16'h00AA;
defparam \saddrInvalid~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Add0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(csr_io_alu_op2_0),
	.datad(csr_io_alu_op1_0),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'h0FF0;
defparam \Add0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Add0~1 (
	.dataa(csr_io_alu_op2_0),
	.datab(csr_io_alu_op1_0),
	.datac(csr_io_alu_op1_1),
	.datad(csr_io_alu_op2_1),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
defparam \Add0~1 .lut_mask = 16'h8778;
defparam \Add0~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \laddrInvalid~1 (
	.dataa(ex_ctrl_mask_type_1),
	.datab(\Add0~0_combout ),
	.datac(\Add0~1_combout ),
	.datad(ex_ctrl_mask_type_0),
	.cin(gnd),
	.combout(\laddrInvalid~1_combout ),
	.cout());
defparam \laddrInvalid~1 .lut_mask = 16'hA888;
defparam \laddrInvalid~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mcause[0]~5 (
	.dataa(waitrequest_reset_override),
	.datab(wait_latency_counter_0),
	.datac(mem_ctrl_mem_wr10),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\mcause[0]~5_combout ),
	.cout());
defparam \mcause[0]~5 .lut_mask = 16'h0028;
defparam \mcause[0]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~0 (
	.dataa(ex_npc_0),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~0_combout ),
	.cout());
defparam \pre_mepc~0 .lut_mask = 16'h8888;
defparam \pre_mepc~0 .sum_lutc_input = "datac";

dffeas \pre_mepc[0] (
	.clk(clock),
	.d(\pre_mepc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[0]~q ),
	.prn(vcc));
defparam \pre_mepc[0] .is_wysiwyg = "true";
defparam \pre_mepc[0] .power_up = "low";

cyclone10lp_lcell_comb \_GEN_204[0]~0 (
	.dataa(\pre_mepc[0]~q ),
	.datab(ex_npc_0),
	.datac(ex_npc_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\_GEN_204[0]~0_combout ),
	.cout());
defparam \_GEN_204[0]~0 .lut_mask = 16'hA8A8;
defparam \_GEN_204[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_246[0]~1 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_0),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_246[0]~1_combout ),
	.cout());
defparam \_T_246[0]~1 .lut_mask = 16'h002A;
defparam \_T_246[0]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_246[0]~2 (
	.dataa(io_out_0),
	.datab(csr_io_in_0),
	.datac(\_T_246[0]~0_combout ),
	.datad(\_T_246[0]~1_combout ),
	.cin(gnd),
	.combout(\_T_246[0]~2_combout ),
	.cout());
defparam \_T_246[0]~2 .lut_mask = 16'hEAC0;
defparam \_T_246[0]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_246[0]~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~0_combout ),
	.cout());
defparam \mtvec~0 .lut_mask = 16'h8888;
defparam \mtvec~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal19~1 (
	.dataa(\Equal19~0_combout ),
	.datab(\Equal16~0_combout ),
	.datac(gnd),
	.datad(ex_csr_addr_11),
	.cin(gnd),
	.combout(\Equal19~1_combout ),
	.cout());
defparam \Equal19~1 .lut_mask = 16'h0088;
defparam \Equal19~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal19~2 (
	.dataa(ex_csr_addr_0),
	.datab(gnd),
	.datac(ex_csr_addr_1),
	.datad(ex_csr_addr_6),
	.cin(gnd),
	.combout(\Equal19~2_combout ),
	.cout());
defparam \Equal19~2 .lut_mask = 16'h000A;
defparam \Equal19~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal19~3 (
	.dataa(ex_csr_addr_2),
	.datab(\Equal19~1_combout ),
	.datac(\Equal19~2_combout ),
	.datad(ex_csr_addr_10),
	.cin(gnd),
	.combout(\Equal19~3_combout ),
	.cout());
defparam \Equal19~3 .lut_mask = 16'h0080;
defparam \Equal19~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \instreth~32 (
	.dataa(io_expt1),
	.datab(mcause_0),
	.datac(\wen~combout ),
	.datad(isEcall),
	.cin(gnd),
	.combout(\instreth~32_combout ),
	.cout());
defparam \instreth~32 .lut_mask = 16'h0080;
defparam \instreth~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec[5]~1 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(gnd),
	.datac(\Equal19~3_combout ),
	.datad(\instreth~32_combout ),
	.cin(gnd),
	.combout(\mtvec[5]~1_combout ),
	.cout());
defparam \mtvec[5]~1 .lut_mask = 16'hF555;
defparam \mtvec[5]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \pre_mepc~2 (
	.dataa(ex_npc_1),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pre_mepc~2_combout ),
	.cout());
defparam \pre_mepc~2 .lut_mask = 16'h8888;
defparam \pre_mepc~2 .sum_lutc_input = "datac";

dffeas \pre_mepc[1] (
	.clk(clock),
	.d(\pre_mepc~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pre_mepc[28]~1_combout ),
	.q(\pre_mepc[1]~q ),
	.prn(vcc));
defparam \pre_mepc[1] .is_wysiwyg = "true";
defparam \pre_mepc[1] .power_up = "low";

cyclone10lp_lcell_comb \_GEN_204[1]~1 (
	.dataa(\pre_mepc[1]~q ),
	.datab(ex_npc_0),
	.datac(ex_npc_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\_GEN_204[1]~1_combout ),
	.cout());
defparam \_GEN_204[1]~1 .lut_mask = 16'hA8A8;
defparam \_GEN_204[1]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_246[1]~3 (
	.dataa(ex_csr_cmd_1),
	.datab(ex_csr_cmd_0),
	.datac(csr_io_in_1),
	.datad(ex_csr_cmd_2),
	.cin(gnd),
	.combout(\_T_246[1]~3_combout ),
	.cout());
defparam \_T_246[1]~3 .lut_mask = 16'h002A;
defparam \_T_246[1]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_246[1]~4 (
	.dataa(io_out_1),
	.datab(\_T_246[0]~0_combout ),
	.datac(csr_io_in_1),
	.datad(\_T_246[1]~3_combout ),
	.cin(gnd),
	.combout(\_T_246[1]~4_combout ),
	.cout());
defparam \_T_246[1]~4 .lut_mask = 16'hEAC0;
defparam \_T_246[1]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_246[1]~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~2_combout ),
	.cout());
defparam \mtvec~2 .lut_mask = 16'h8888;
defparam \mtvec~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal30~0 (
	.dataa(Equal62),
	.datab(\Equal25~2_combout ),
	.datac(\Equal16~0_combout ),
	.datad(ex_csr_addr_6),
	.cin(gnd),
	.combout(\Equal30~0_combout ),
	.cout());
defparam \Equal30~0 .lut_mask = 16'h0080;
defparam \Equal30~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal25~3 (
	.dataa(Equal62),
	.datab(ex_csr_addr_6),
	.datac(\Equal25~2_combout ),
	.datad(\Equal16~0_combout ),
	.cin(gnd),
	.combout(\Equal25~3_combout ),
	.cout());
defparam \Equal25~3 .lut_mask = 16'h8000;
defparam \Equal25~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mscratch[0]~0 (
	.dataa(\Equal25~3_combout ),
	.datab(\instreth~32_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mscratch[0]~0_combout ),
	.cout());
defparam \mscratch[0]~0 .lut_mask = 16'h8888;
defparam \mscratch[0]~0 .sum_lutc_input = "datac";

dffeas \mscratch[1] (
	.clk(clock),
	.d(\_T_246[1]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[1]~q ),
	.prn(vcc));
defparam \mscratch[1] .is_wysiwyg = "true";
defparam \mscratch[1] .power_up = "low";

cyclone10lp_lcell_comb \io_out[1]~2 (
	.dataa(\Equal30~0_combout ),
	.datab(\Equal25~3_combout ),
	.datac(\mscratch[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[1]~2_combout ),
	.cout());
defparam \io_out[1]~2 .lut_mask = 16'hEAEA;
defparam \io_out[1]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal16~1 (
	.dataa(\Equal19~0_combout ),
	.datab(ex_csr_addr_11),
	.datac(ex_csr_addr_2),
	.datad(ex_csr_addr_6),
	.cin(gnd),
	.combout(\Equal16~1_combout ),
	.cout());
defparam \Equal16~1 .lut_mask = 16'h0008;
defparam \Equal16~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal3~0 (
	.dataa(ex_csr_addr_10),
	.datab(\Equal16~1_combout ),
	.datac(ex_csr_addr_8),
	.datad(ex_csr_addr_9),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
defparam \Equal3~0 .lut_mask = 16'h0008;
defparam \Equal3~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal11~2 (
	.dataa(ex_csr_addr_8),
	.datab(\Equal16~1_combout ),
	.datac(ex_csr_addr_10),
	.datad(ex_csr_addr_9),
	.cin(gnd),
	.combout(\Equal11~2_combout ),
	.cout());
defparam \Equal11~2 .lut_mask = 16'h0008;
defparam \Equal11~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal11~3 (
	.dataa(ex_csr_addr_0),
	.datab(ex_csr_addr_1),
	.datac(\Equal11~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal11~3_combout ),
	.cout());
defparam \Equal11~3 .lut_mask = 16'h2020;
defparam \Equal11~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal23~0 (
	.dataa(ex_csr_addr_10),
	.datab(\Equal4~0_combout ),
	.datac(\Equal19~1_combout ),
	.datad(ex_csr_addr_2),
	.cin(gnd),
	.combout(\Equal23~0_combout ),
	.cout());
defparam \Equal23~0 .lut_mask = 16'h0080;
defparam \Equal23~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[1]~3 (
	.dataa(ex_csr_addr_6),
	.datab(ex_csr_addr_7),
	.datac(\Equal11~3_combout ),
	.datad(\Equal23~0_combout ),
	.cin(gnd),
	.combout(\io_out[1]~3_combout ),
	.cout());
defparam \io_out[1]~3 .lut_mask = 16'h8ACF;
defparam \io_out[1]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[1]~4 (
	.dataa(\Equal4~0_combout ),
	.datab(\Equal3~0_combout ),
	.datac(ex_csr_addr_7),
	.datad(\io_out[1]~3_combout ),
	.cin(gnd),
	.combout(\io_out[1]~4_combout ),
	.cout());
defparam \io_out[1]~4 .lut_mask = 16'h08FF;
defparam \io_out[1]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \time_[0]~32 (
	.dataa(\time_[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\time_[0]~32_combout ),
	.cout(\time_[0]~33 ));
defparam \time_[0]~32 .lut_mask = 16'h55AA;
defparam \time_[0]~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal19~4 (
	.dataa(ex_csr_addr_2),
	.datab(\Equal19~1_combout ),
	.datac(gnd),
	.datad(ex_csr_addr_10),
	.cin(gnd),
	.combout(\Equal19~4_combout ),
	.cout());
defparam \Equal19~4 .lut_mask = 16'h0088;
defparam \Equal19~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal21~2 (
	.dataa(ex_csr_addr_0),
	.datab(ex_csr_addr_1),
	.datac(\Equal19~4_combout ),
	.datad(ex_csr_addr_6),
	.cin(gnd),
	.combout(\Equal21~2_combout ),
	.cout());
defparam \Equal21~2 .lut_mask = 16'h0010;
defparam \Equal21~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal29~2 (
	.dataa(ex_csr_addr_0),
	.datab(ex_csr_addr_1),
	.datac(ex_csr_addr_6),
	.datad(\Equal19~4_combout ),
	.cin(gnd),
	.combout(\Equal29~2_combout ),
	.cout());
defparam \Equal29~2 .lut_mask = 16'h1000;
defparam \Equal29~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \timeh~33 (
	.dataa(\instreth~32_combout ),
	.datab(\Equal30~0_combout ),
	.datac(\Equal21~2_combout ),
	.datad(\Equal29~2_combout ),
	.cin(gnd),
	.combout(\timeh~33_combout ),
	.cout());
defparam \timeh~33 .lut_mask = 16'h0002;
defparam \timeh~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \time_~36 (
	.dataa(\timeh~33_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\io_out[1]~3_combout ),
	.cin(gnd),
	.combout(\time_~36_combout ),
	.cout());
defparam \time_~36 .lut_mask = 16'h00AA;
defparam \time_~36 .sum_lutc_input = "datac";

dffeas \time_[0] (
	.clk(clock),
	.d(\time_[0]~32_combout ),
	.asdata(\_T_246[0]~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[0]~q ),
	.prn(vcc));
defparam \time_[0] .is_wysiwyg = "true";
defparam \time_[0] .power_up = "low";

cyclone10lp_lcell_comb \time_[1]~34 (
	.dataa(\time_[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[0]~33 ),
	.combout(\time_[1]~34_combout ),
	.cout(\time_[1]~35 ));
defparam \time_[1]~34 .lut_mask = 16'h5A5F;
defparam \time_[1]~34 .sum_lutc_input = "cin";

dffeas \time_[1] (
	.clk(clock),
	.d(\time_[1]~34_combout ),
	.asdata(\_T_246[1]~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[1]~q ),
	.prn(vcc));
defparam \time_[1] .is_wysiwyg = "true";
defparam \time_[1] .power_up = "low";

cyclone10lp_lcell_comb \io_out[1]~5 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_1),
	.datad(\time_[1]~q ),
	.cin(gnd),
	.combout(\io_out[1]~5_combout ),
	.cout());
defparam \io_out[1]~5 .lut_mask = 16'hEAC0;
defparam \io_out[1]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal9~0 (
	.dataa(\Equal11~2_combout ),
	.datab(ex_csr_addr_0),
	.datac(ex_csr_addr_1),
	.datad(ex_csr_addr_7),
	.cin(gnd),
	.combout(\Equal9~0_combout ),
	.cout());
defparam \Equal9~0 .lut_mask = 16'h0002;
defparam \Equal9~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[1]~6 (
	.dataa(\Equal9~0_combout ),
	.datab(Equal62),
	.datac(\Equal3~0_combout ),
	.datad(ex_csr_addr_7),
	.cin(gnd),
	.combout(\io_out[1]~6_combout ),
	.cout());
defparam \io_out[1]~6 .lut_mask = 16'hAAEA;
defparam \io_out[1]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cycle[0]~32 (
	.dataa(\cycle[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\cycle[0]~32_combout ),
	.cout(\cycle[0]~33 ));
defparam \cycle[0]~32 .lut_mask = 16'h55AA;
defparam \cycle[0]~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cycle~36 (
	.dataa(\Equal9~0_combout ),
	.datab(\instreth~32_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\cycle~36_combout ),
	.cout());
defparam \cycle~36 .lut_mask = 16'h8888;
defparam \cycle~36 .sum_lutc_input = "datac";

dffeas \cycle[0] (
	.clk(clock),
	.d(\cycle[0]~32_combout ),
	.asdata(\_T_246[0]~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[0]~q ),
	.prn(vcc));
defparam \cycle[0] .is_wysiwyg = "true";
defparam \cycle[0] .power_up = "low";

cyclone10lp_lcell_comb \cycle[1]~34 (
	.dataa(\cycle[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[0]~33 ),
	.combout(\cycle[1]~34_combout ),
	.cout(\cycle[1]~35 ));
defparam \cycle[1]~34 .lut_mask = 16'h5A5F;
defparam \cycle[1]~34 .sum_lutc_input = "cin";

dffeas \cycle[1] (
	.clk(clock),
	.d(\cycle[1]~34_combout ),
	.asdata(\_T_246[1]~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[1]~q ),
	.prn(vcc));
defparam \cycle[1] .is_wysiwyg = "true";
defparam \cycle[1] .power_up = "low";

cyclone10lp_lcell_comb \io_out[1]~7 (
	.dataa(\io_out[1]~2_combout ),
	.datab(\io_out[1]~5_combout ),
	.datac(\io_out[1]~6_combout ),
	.datad(\cycle[1]~q ),
	.cin(gnd),
	.combout(\io_out[1]~7_combout ),
	.cout());
defparam \io_out[1]~7 .lut_mask = 16'hFEEE;
defparam \io_out[1]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal25~5 (
	.dataa(ex_csr_addr_8),
	.datab(ex_csr_addr_9),
	.datac(ex_csr_addr_7),
	.datad(\Equal25~2_combout ),
	.cin(gnd),
	.combout(\Equal25~5_combout ),
	.cout());
defparam \Equal25~5 .lut_mask = 16'h0800;
defparam \Equal25~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal27~0 (
	.dataa(ex_csr_addr_1),
	.datab(ex_csr_addr_6),
	.datac(\Equal25~5_combout ),
	.datad(ex_csr_addr_0),
	.cin(gnd),
	.combout(\Equal27~0_combout ),
	.cout());
defparam \Equal27~0 .lut_mask = 16'h0080;
defparam \Equal27~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal12~0 (
	.dataa(ex_csr_addr_1),
	.datab(\Equal11~2_combout ),
	.datac(ex_csr_addr_0),
	.datad(ex_csr_addr_7),
	.cin(gnd),
	.combout(\Equal12~0_combout ),
	.cout());
defparam \Equal12~0 .lut_mask = 16'h0008;
defparam \Equal12~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal8~0 (
	.dataa(ex_csr_addr_1),
	.datab(\Equal3~0_combout ),
	.datac(gnd),
	.datad(ex_csr_addr_0),
	.cin(gnd),
	.combout(\Equal8~0_combout ),
	.cout());
defparam \Equal8~0 .lut_mask = 16'h0088;
defparam \Equal8~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[1]~8 (
	.dataa(\Equal12~0_combout ),
	.datab(\Equal8~0_combout ),
	.datac(gnd),
	.datad(ex_csr_addr_7),
	.cin(gnd),
	.combout(\io_out[1]~8_combout ),
	.cout());
defparam \io_out[1]~8 .lut_mask = 16'hAAEE;
defparam \io_out[1]~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \instret[0]~34 (
	.dataa(\instret[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\instret[0]~34_combout ),
	.cout(\instret[0]~35 ));
defparam \instret[0]~34 .lut_mask = 16'h55AA;
defparam \instret[0]~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \instret~38 (
	.dataa(\Equal12~0_combout ),
	.datab(\instreth~32_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instret~38_combout ),
	.cout());
defparam \instret~38 .lut_mask = 16'h8888;
defparam \instret~38 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal39~0 (
	.dataa(ex_csr_addr_0),
	.datab(ex_csr_addr_1),
	.datac(ex_csr_addr_6),
	.datad(ex_csr_addr_7),
	.cin(gnd),
	.combout(\Equal39~0_combout ),
	.cout());
defparam \Equal39~0 .lut_mask = 16'h0001;
defparam \Equal39~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal39~1 (
	.dataa(ex_inst_0),
	.datab(ex_inst_1),
	.datac(ex_csr_addr_8),
	.datad(ex_csr_addr_9),
	.cin(gnd),
	.combout(\Equal39~1_combout ),
	.cout());
defparam \Equal39~1 .lut_mask = 16'h0008;
defparam \Equal39~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal39~2 (
	.dataa(ex_inst_4),
	.datab(ex_inst_2),
	.datac(ex_inst_3),
	.datad(ex_inst_5),
	.cin(gnd),
	.combout(\Equal39~2_combout ),
	.cout());
defparam \Equal39~2 .lut_mask = 16'h0002;
defparam \Equal39~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal39~3 (
	.dataa(ex_inst_7),
	.datab(ex_inst_8),
	.datac(ex_inst_9),
	.datad(ex_inst_6),
	.cin(gnd),
	.combout(\Equal39~3_combout ),
	.cout());
defparam \Equal39~3 .lut_mask = 16'h0001;
defparam \Equal39~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal39~4 (
	.dataa(\Equal39~0_combout ),
	.datab(\Equal39~1_combout ),
	.datac(\Equal39~2_combout ),
	.datad(\Equal39~3_combout ),
	.cin(gnd),
	.combout(\Equal39~4_combout ),
	.cout());
defparam \Equal39~4 .lut_mask = 16'h8000;
defparam \Equal39~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal39~5 (
	.dataa(ex_inst_11),
	.datab(ex_inst_10),
	.datac(ex_inst_12),
	.datad(ex_inst_13),
	.cin(gnd),
	.combout(\Equal39~5_combout ),
	.cout());
defparam \Equal39~5 .lut_mask = 16'h0001;
defparam \Equal39~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal39~6 (
	.dataa(\Equal39~4_combout ),
	.datab(\Equal39~5_combout ),
	.datac(gnd),
	.datad(ex_inst_14),
	.cin(gnd),
	.combout(\Equal39~6_combout ),
	.cout());
defparam \Equal39~6 .lut_mask = 16'h0088;
defparam \Equal39~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \isInstRet~0 (
	.dataa(Equal59),
	.datab(\Equal25~2_combout ),
	.datac(\Equal39~6_combout ),
	.datad(mcause_0),
	.cin(gnd),
	.combout(\isInstRet~0_combout ),
	.cout());
defparam \isInstRet~0 .lut_mask = 16'h80FF;
defparam \isInstRet~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \instret[0]~99 (
	.dataa(\isInstRet~0_combout ),
	.datab(io_expt1),
	.datac(isEcall),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\instret[0]~99_combout ),
	.cout());
defparam \instret[0]~99 .lut_mask = 16'h54FF;
defparam \instret[0]~99 .sum_lutc_input = "datac";

dffeas \instret[0] (
	.clk(clock),
	.d(\instret[0]~34_combout ),
	.asdata(\_T_246[0]~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[0]~q ),
	.prn(vcc));
defparam \instret[0] .is_wysiwyg = "true";
defparam \instret[0] .power_up = "low";

cyclone10lp_lcell_comb \instret[1]~36 (
	.dataa(\instret[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[0]~35 ),
	.combout(\instret[1]~36_combout ),
	.cout(\instret[1]~37 ));
defparam \instret[1]~36 .lut_mask = 16'h5A5F;
defparam \instret[1]~36 .sum_lutc_input = "cin";

dffeas \instret[1] (
	.clk(clock),
	.d(\instret[1]~36_combout ),
	.asdata(\_T_246[1]~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[1]~q ),
	.prn(vcc));
defparam \instret[1] .is_wysiwyg = "true";
defparam \instret[1] .power_up = "low";

cyclone10lp_lcell_comb \mcause[2]~7 (
	.dataa(\mcause~4_combout ),
	.datab(\laddrInvalid~0_combout ),
	.datac(\laddrInvalid~1_combout ),
	.datad(isEcall),
	.cin(gnd),
	.combout(\mcause[2]~7_combout ),
	.cout());
defparam \mcause[2]~7 .lut_mask = 16'h008A;
defparam \mcause[2]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_219~0 (
	.dataa(Equal56),
	.datab(\Add0~0_combout ),
	.datac(\Add0~1_combout ),
	.datad(ex_j_check),
	.cin(gnd),
	.combout(\_T_219~0_combout ),
	.cout());
defparam \_T_219~0 .lut_mask = 16'h02AA;
defparam \_T_219~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mcause~8 (
	.dataa(\mcause[2]~7_combout ),
	.datab(\_T_219~0_combout ),
	.datac(\isIllegal~0_combout ),
	.datad(isEcall),
	.cin(gnd),
	.combout(\mcause~8_combout ),
	.cout());
defparam \mcause~8 .lut_mask = 16'hFFAE;
defparam \mcause~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \saddrInvalid~1 (
	.dataa(ex_ctrl_imm_type001),
	.datab(\laddrInvalid~1_combout ),
	.datac(gnd),
	.datad(ex_ctrl_mask_type_2),
	.cin(gnd),
	.combout(\saddrInvalid~1_combout ),
	.cout());
defparam \saddrInvalid~1 .lut_mask = 16'h0088;
defparam \saddrInvalid~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mcause~9 (
	.dataa(\saddrInvalid~1_combout ),
	.datab(isEcall),
	.datac(io_expt1),
	.datad(\mcause[2]~7_combout ),
	.cin(gnd),
	.combout(\mcause~9_combout ),
	.cout());
defparam \mcause~9 .lut_mask = 16'h8ACF;
defparam \mcause~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mcause~10 (
	.dataa(io_expt2),
	.datab(\mcause~8_combout ),
	.datac(\mcause~9_combout ),
	.datad(\_T_246[1]~4_combout ),
	.cin(gnd),
	.combout(\mcause~10_combout ),
	.cout());
defparam \mcause~10 .lut_mask = 16'hEAC0;
defparam \mcause~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mcause[0]~11 (
	.dataa(mcause_0),
	.datab(\Equal27~0_combout ),
	.datac(\wen~combout ),
	.datad(io_expt2),
	.cin(gnd),
	.combout(\mcause[0]~11_combout ),
	.cout());
defparam \mcause[0]~11 .lut_mask = 16'h80AA;
defparam \mcause[0]~11 .sum_lutc_input = "datac";

dffeas \mcause[1] (
	.clk(clock),
	.d(\mcause~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mcause[0]~11_combout ),
	.q(\mcause[1]~q ),
	.prn(vcc));
defparam \mcause[1] .is_wysiwyg = "true";
defparam \mcause[1] .power_up = "low";

cyclone10lp_lcell_comb \io_out[1]~9 (
	.dataa(\Equal27~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[1]~q ),
	.datad(\mcause[1]~q ),
	.cin(gnd),
	.combout(\io_out[1]~9_combout ),
	.cout());
defparam \io_out[1]~9 .lut_mask = 16'hEAC0;
defparam \io_out[1]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal28~0 (
	.dataa(ex_csr_addr_0),
	.datab(ex_csr_addr_1),
	.datac(ex_csr_addr_6),
	.datad(\Equal25~5_combout ),
	.cin(gnd),
	.combout(\Equal28~0_combout ),
	.cout());
defparam \Equal28~0 .lut_mask = 16'h8000;
defparam \Equal28~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal13~0 (
	.dataa(ex_csr_addr_7),
	.datab(\Equal11~2_combout ),
	.datac(ex_csr_addr_0),
	.datad(ex_csr_addr_1),
	.cin(gnd),
	.combout(\Equal13~0_combout ),
	.cout());
defparam \Equal13~0 .lut_mask = 16'h0008;
defparam \Equal13~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[1]~10 (
	.dataa(\Equal13~0_combout ),
	.datab(Equal62),
	.datac(ex_csr_addr_7),
	.datad(\Equal3~0_combout ),
	.cin(gnd),
	.combout(\io_out[1]~10_combout ),
	.cout());
defparam \io_out[1]~10 .lut_mask = 16'hEAAA;
defparam \io_out[1]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cycleh[0]~32 (
	.dataa(\cycleh[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\cycleh[0]~32_combout ),
	.cout(\cycleh[0]~33 ));
defparam \cycleh[0]~32 .lut_mask = 16'h55AA;
defparam \cycleh[0]~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cycleh~36 (
	.dataa(\Equal13~0_combout ),
	.datab(\instreth~32_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\cycleh~36_combout ),
	.cout());
defparam \cycleh~36 .lut_mask = 16'h8888;
defparam \cycleh~36 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cycle[2]~37 (
	.dataa(\cycle[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[1]~35 ),
	.combout(\cycle[2]~37_combout ),
	.cout(\cycle[2]~38 ));
defparam \cycle[2]~37 .lut_mask = 16'hA50A;
defparam \cycle[2]~37 .sum_lutc_input = "cin";

dffeas \cycle[2] (
	.clk(clock),
	.d(\cycle[2]~37_combout ),
	.asdata(\_T_246[2]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[2]~q ),
	.prn(vcc));
defparam \cycle[2] .is_wysiwyg = "true";
defparam \cycle[2] .power_up = "low";

cyclone10lp_lcell_comb \cycle[3]~39 (
	.dataa(\cycle[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[2]~38 ),
	.combout(\cycle[3]~39_combout ),
	.cout(\cycle[3]~40 ));
defparam \cycle[3]~39 .lut_mask = 16'h5A5F;
defparam \cycle[3]~39 .sum_lutc_input = "cin";

dffeas \cycle[3] (
	.clk(clock),
	.d(\cycle[3]~39_combout ),
	.asdata(\_T_246[3]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[3]~q ),
	.prn(vcc));
defparam \cycle[3] .is_wysiwyg = "true";
defparam \cycle[3] .power_up = "low";

cyclone10lp_lcell_comb \cycle[4]~41 (
	.dataa(\cycle[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[3]~40 ),
	.combout(\cycle[4]~41_combout ),
	.cout(\cycle[4]~42 ));
defparam \cycle[4]~41 .lut_mask = 16'hA50A;
defparam \cycle[4]~41 .sum_lutc_input = "cin";

dffeas \cycle[4] (
	.clk(clock),
	.d(\cycle[4]~41_combout ),
	.asdata(\_T_244[4]~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[4]~q ),
	.prn(vcc));
defparam \cycle[4] .is_wysiwyg = "true";
defparam \cycle[4] .power_up = "low";

cyclone10lp_lcell_comb \cycle[5]~43 (
	.dataa(\cycle[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[4]~42 ),
	.combout(\cycle[5]~43_combout ),
	.cout(\cycle[5]~44 ));
defparam \cycle[5]~43 .lut_mask = 16'h5A5F;
defparam \cycle[5]~43 .sum_lutc_input = "cin";

dffeas \cycle[5] (
	.clk(clock),
	.d(\cycle[5]~43_combout ),
	.asdata(\_T_244[5]~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[5]~q ),
	.prn(vcc));
defparam \cycle[5] .is_wysiwyg = "true";
defparam \cycle[5] .power_up = "low";

cyclone10lp_lcell_comb \cycle[6]~45 (
	.dataa(\cycle[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[5]~44 ),
	.combout(\cycle[6]~45_combout ),
	.cout(\cycle[6]~46 ));
defparam \cycle[6]~45 .lut_mask = 16'hA50A;
defparam \cycle[6]~45 .sum_lutc_input = "cin";

dffeas \cycle[6] (
	.clk(clock),
	.d(\cycle[6]~45_combout ),
	.asdata(\_T_244[6]~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[6]~q ),
	.prn(vcc));
defparam \cycle[6] .is_wysiwyg = "true";
defparam \cycle[6] .power_up = "low";

cyclone10lp_lcell_comb \cycle[7]~47 (
	.dataa(\cycle[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[6]~46 ),
	.combout(\cycle[7]~47_combout ),
	.cout(\cycle[7]~48 ));
defparam \cycle[7]~47 .lut_mask = 16'h5A5F;
defparam \cycle[7]~47 .sum_lutc_input = "cin";

dffeas \cycle[7] (
	.clk(clock),
	.d(\cycle[7]~47_combout ),
	.asdata(\_T_244[7]~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[7]~q ),
	.prn(vcc));
defparam \cycle[7] .is_wysiwyg = "true";
defparam \cycle[7] .power_up = "low";

cyclone10lp_lcell_comb \cycle[8]~49 (
	.dataa(\cycle[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[7]~48 ),
	.combout(\cycle[8]~49_combout ),
	.cout(\cycle[8]~50 ));
defparam \cycle[8]~49 .lut_mask = 16'hA50A;
defparam \cycle[8]~49 .sum_lutc_input = "cin";

dffeas \cycle[8] (
	.clk(clock),
	.d(\cycle[8]~49_combout ),
	.asdata(\_T_244[8]~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[8]~q ),
	.prn(vcc));
defparam \cycle[8] .is_wysiwyg = "true";
defparam \cycle[8] .power_up = "low";

cyclone10lp_lcell_comb \cycle[9]~51 (
	.dataa(\cycle[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[8]~50 ),
	.combout(\cycle[9]~51_combout ),
	.cout(\cycle[9]~52 ));
defparam \cycle[9]~51 .lut_mask = 16'h5A5F;
defparam \cycle[9]~51 .sum_lutc_input = "cin";

dffeas \cycle[9] (
	.clk(clock),
	.d(\cycle[9]~51_combout ),
	.asdata(\_T_244[9]~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[9]~q ),
	.prn(vcc));
defparam \cycle[9] .is_wysiwyg = "true";
defparam \cycle[9] .power_up = "low";

cyclone10lp_lcell_comb \cycle[10]~53 (
	.dataa(\cycle[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[9]~52 ),
	.combout(\cycle[10]~53_combout ),
	.cout(\cycle[10]~54 ));
defparam \cycle[10]~53 .lut_mask = 16'hA50A;
defparam \cycle[10]~53 .sum_lutc_input = "cin";

dffeas \cycle[10] (
	.clk(clock),
	.d(\cycle[10]~53_combout ),
	.asdata(\_T_244[10]~13_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[10]~q ),
	.prn(vcc));
defparam \cycle[10] .is_wysiwyg = "true";
defparam \cycle[10] .power_up = "low";

cyclone10lp_lcell_comb \cycle[11]~55 (
	.dataa(\cycle[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[10]~54 ),
	.combout(\cycle[11]~55_combout ),
	.cout(\cycle[11]~56 ));
defparam \cycle[11]~55 .lut_mask = 16'h5A5F;
defparam \cycle[11]~55 .sum_lutc_input = "cin";

dffeas \cycle[11] (
	.clk(clock),
	.d(\cycle[11]~55_combout ),
	.asdata(\_T_244[11]~15_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[11]~q ),
	.prn(vcc));
defparam \cycle[11] .is_wysiwyg = "true";
defparam \cycle[11] .power_up = "low";

cyclone10lp_lcell_comb \cycle[12]~57 (
	.dataa(\cycle[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[11]~56 ),
	.combout(\cycle[12]~57_combout ),
	.cout(\cycle[12]~58 ));
defparam \cycle[12]~57 .lut_mask = 16'hA50A;
defparam \cycle[12]~57 .sum_lutc_input = "cin";

dffeas \cycle[12] (
	.clk(clock),
	.d(\cycle[12]~57_combout ),
	.asdata(\_T_244[12]~17_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[12]~q ),
	.prn(vcc));
defparam \cycle[12] .is_wysiwyg = "true";
defparam \cycle[12] .power_up = "low";

cyclone10lp_lcell_comb \cycle[13]~59 (
	.dataa(\cycle[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[12]~58 ),
	.combout(\cycle[13]~59_combout ),
	.cout(\cycle[13]~60 ));
defparam \cycle[13]~59 .lut_mask = 16'h5A5F;
defparam \cycle[13]~59 .sum_lutc_input = "cin";

dffeas \cycle[13] (
	.clk(clock),
	.d(\cycle[13]~59_combout ),
	.asdata(\_T_244[13]~19_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[13]~q ),
	.prn(vcc));
defparam \cycle[13] .is_wysiwyg = "true";
defparam \cycle[13] .power_up = "low";

cyclone10lp_lcell_comb \cycle[14]~61 (
	.dataa(\cycle[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[13]~60 ),
	.combout(\cycle[14]~61_combout ),
	.cout(\cycle[14]~62 ));
defparam \cycle[14]~61 .lut_mask = 16'hA50A;
defparam \cycle[14]~61 .sum_lutc_input = "cin";

dffeas \cycle[14] (
	.clk(clock),
	.d(\cycle[14]~61_combout ),
	.asdata(\_T_244[14]~21_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[14]~q ),
	.prn(vcc));
defparam \cycle[14] .is_wysiwyg = "true";
defparam \cycle[14] .power_up = "low";

cyclone10lp_lcell_comb \cycle[15]~63 (
	.dataa(\cycle[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[14]~62 ),
	.combout(\cycle[15]~63_combout ),
	.cout(\cycle[15]~64 ));
defparam \cycle[15]~63 .lut_mask = 16'h5A5F;
defparam \cycle[15]~63 .sum_lutc_input = "cin";

dffeas \cycle[15] (
	.clk(clock),
	.d(\cycle[15]~63_combout ),
	.asdata(\_T_244[15]~23_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[15]~q ),
	.prn(vcc));
defparam \cycle[15] .is_wysiwyg = "true";
defparam \cycle[15] .power_up = "low";

cyclone10lp_lcell_comb \cycle[16]~65 (
	.dataa(\cycle[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[15]~64 ),
	.combout(\cycle[16]~65_combout ),
	.cout(\cycle[16]~66 ));
defparam \cycle[16]~65 .lut_mask = 16'hA50A;
defparam \cycle[16]~65 .sum_lutc_input = "cin";

dffeas \cycle[16] (
	.clk(clock),
	.d(\cycle[16]~65_combout ),
	.asdata(\_T_244[16]~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[16]~q ),
	.prn(vcc));
defparam \cycle[16] .is_wysiwyg = "true";
defparam \cycle[16] .power_up = "low";

cyclone10lp_lcell_comb \cycle[17]~67 (
	.dataa(\cycle[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[16]~66 ),
	.combout(\cycle[17]~67_combout ),
	.cout(\cycle[17]~68 ));
defparam \cycle[17]~67 .lut_mask = 16'h5A5F;
defparam \cycle[17]~67 .sum_lutc_input = "cin";

dffeas \cycle[17] (
	.clk(clock),
	.d(\cycle[17]~67_combout ),
	.asdata(\_T_244[17]~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[17]~q ),
	.prn(vcc));
defparam \cycle[17] .is_wysiwyg = "true";
defparam \cycle[17] .power_up = "low";

cyclone10lp_lcell_comb \cycle[18]~69 (
	.dataa(\cycle[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[17]~68 ),
	.combout(\cycle[18]~69_combout ),
	.cout(\cycle[18]~70 ));
defparam \cycle[18]~69 .lut_mask = 16'hA50A;
defparam \cycle[18]~69 .sum_lutc_input = "cin";

dffeas \cycle[18] (
	.clk(clock),
	.d(\cycle[18]~69_combout ),
	.asdata(\_T_244[18]~29_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[18]~q ),
	.prn(vcc));
defparam \cycle[18] .is_wysiwyg = "true";
defparam \cycle[18] .power_up = "low";

cyclone10lp_lcell_comb \cycle[19]~71 (
	.dataa(\cycle[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[18]~70 ),
	.combout(\cycle[19]~71_combout ),
	.cout(\cycle[19]~72 ));
defparam \cycle[19]~71 .lut_mask = 16'h5A5F;
defparam \cycle[19]~71 .sum_lutc_input = "cin";

dffeas \cycle[19] (
	.clk(clock),
	.d(\cycle[19]~71_combout ),
	.asdata(\_T_244[19]~31_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[19]~q ),
	.prn(vcc));
defparam \cycle[19] .is_wysiwyg = "true";
defparam \cycle[19] .power_up = "low";

cyclone10lp_lcell_comb \cycle[20]~73 (
	.dataa(\cycle[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[19]~72 ),
	.combout(\cycle[20]~73_combout ),
	.cout(\cycle[20]~74 ));
defparam \cycle[20]~73 .lut_mask = 16'hA50A;
defparam \cycle[20]~73 .sum_lutc_input = "cin";

dffeas \cycle[20] (
	.clk(clock),
	.d(\cycle[20]~73_combout ),
	.asdata(\_T_244[20]~33_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[20]~q ),
	.prn(vcc));
defparam \cycle[20] .is_wysiwyg = "true";
defparam \cycle[20] .power_up = "low";

cyclone10lp_lcell_comb \cycle[21]~75 (
	.dataa(\cycle[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[20]~74 ),
	.combout(\cycle[21]~75_combout ),
	.cout(\cycle[21]~76 ));
defparam \cycle[21]~75 .lut_mask = 16'h5A5F;
defparam \cycle[21]~75 .sum_lutc_input = "cin";

dffeas \cycle[21] (
	.clk(clock),
	.d(\cycle[21]~75_combout ),
	.asdata(\_T_244[21]~35_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[21]~q ),
	.prn(vcc));
defparam \cycle[21] .is_wysiwyg = "true";
defparam \cycle[21] .power_up = "low";

cyclone10lp_lcell_comb \cycle[22]~77 (
	.dataa(\cycle[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[21]~76 ),
	.combout(\cycle[22]~77_combout ),
	.cout(\cycle[22]~78 ));
defparam \cycle[22]~77 .lut_mask = 16'hA50A;
defparam \cycle[22]~77 .sum_lutc_input = "cin";

dffeas \cycle[22] (
	.clk(clock),
	.d(\cycle[22]~77_combout ),
	.asdata(\_T_244[22]~37_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[22]~q ),
	.prn(vcc));
defparam \cycle[22] .is_wysiwyg = "true";
defparam \cycle[22] .power_up = "low";

cyclone10lp_lcell_comb \cycle[23]~79 (
	.dataa(\cycle[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[22]~78 ),
	.combout(\cycle[23]~79_combout ),
	.cout(\cycle[23]~80 ));
defparam \cycle[23]~79 .lut_mask = 16'h5A5F;
defparam \cycle[23]~79 .sum_lutc_input = "cin";

dffeas \cycle[23] (
	.clk(clock),
	.d(\cycle[23]~79_combout ),
	.asdata(\_T_244[23]~39_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[23]~q ),
	.prn(vcc));
defparam \cycle[23] .is_wysiwyg = "true";
defparam \cycle[23] .power_up = "low";

cyclone10lp_lcell_comb \cycle[24]~81 (
	.dataa(\cycle[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[23]~80 ),
	.combout(\cycle[24]~81_combout ),
	.cout(\cycle[24]~82 ));
defparam \cycle[24]~81 .lut_mask = 16'hA50A;
defparam \cycle[24]~81 .sum_lutc_input = "cin";

dffeas \cycle[24] (
	.clk(clock),
	.d(\cycle[24]~81_combout ),
	.asdata(\_T_244[24]~41_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[24]~q ),
	.prn(vcc));
defparam \cycle[24] .is_wysiwyg = "true";
defparam \cycle[24] .power_up = "low";

cyclone10lp_lcell_comb \cycle[25]~83 (
	.dataa(\cycle[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[24]~82 ),
	.combout(\cycle[25]~83_combout ),
	.cout(\cycle[25]~84 ));
defparam \cycle[25]~83 .lut_mask = 16'h5A5F;
defparam \cycle[25]~83 .sum_lutc_input = "cin";

dffeas \cycle[25] (
	.clk(clock),
	.d(\cycle[25]~83_combout ),
	.asdata(\_T_244[25]~43_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[25]~q ),
	.prn(vcc));
defparam \cycle[25] .is_wysiwyg = "true";
defparam \cycle[25] .power_up = "low";

cyclone10lp_lcell_comb \cycle[26]~85 (
	.dataa(\cycle[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[25]~84 ),
	.combout(\cycle[26]~85_combout ),
	.cout(\cycle[26]~86 ));
defparam \cycle[26]~85 .lut_mask = 16'hA50A;
defparam \cycle[26]~85 .sum_lutc_input = "cin";

dffeas \cycle[26] (
	.clk(clock),
	.d(\cycle[26]~85_combout ),
	.asdata(\_T_244[26]~45_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[26]~q ),
	.prn(vcc));
defparam \cycle[26] .is_wysiwyg = "true";
defparam \cycle[26] .power_up = "low";

cyclone10lp_lcell_comb \cycle[27]~87 (
	.dataa(\cycle[27]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[26]~86 ),
	.combout(\cycle[27]~87_combout ),
	.cout(\cycle[27]~88 ));
defparam \cycle[27]~87 .lut_mask = 16'h5A5F;
defparam \cycle[27]~87 .sum_lutc_input = "cin";

dffeas \cycle[27] (
	.clk(clock),
	.d(\cycle[27]~87_combout ),
	.asdata(\_T_244[27]~47_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[27]~q ),
	.prn(vcc));
defparam \cycle[27] .is_wysiwyg = "true";
defparam \cycle[27] .power_up = "low";

cyclone10lp_lcell_comb \cycle[28]~89 (
	.dataa(\cycle[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[27]~88 ),
	.combout(\cycle[28]~89_combout ),
	.cout(\cycle[28]~90 ));
defparam \cycle[28]~89 .lut_mask = 16'hA50A;
defparam \cycle[28]~89 .sum_lutc_input = "cin";

dffeas \cycle[28] (
	.clk(clock),
	.d(\cycle[28]~89_combout ),
	.asdata(\_T_244[28]~49_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[28]~q ),
	.prn(vcc));
defparam \cycle[28] .is_wysiwyg = "true";
defparam \cycle[28] .power_up = "low";

cyclone10lp_lcell_comb \cycle[29]~91 (
	.dataa(\cycle[29]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[28]~90 ),
	.combout(\cycle[29]~91_combout ),
	.cout(\cycle[29]~92 ));
defparam \cycle[29]~91 .lut_mask = 16'h5A5F;
defparam \cycle[29]~91 .sum_lutc_input = "cin";

dffeas \cycle[29] (
	.clk(clock),
	.d(\cycle[29]~91_combout ),
	.asdata(\_T_244[29]~51_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[29]~q ),
	.prn(vcc));
defparam \cycle[29] .is_wysiwyg = "true";
defparam \cycle[29] .power_up = "low";

cyclone10lp_lcell_comb \cycle[30]~93 (
	.dataa(\cycle[30]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycle[29]~92 ),
	.combout(\cycle[30]~93_combout ),
	.cout(\cycle[30]~94 ));
defparam \cycle[30]~93 .lut_mask = 16'hA50A;
defparam \cycle[30]~93 .sum_lutc_input = "cin";

dffeas \cycle[30] (
	.clk(clock),
	.d(\cycle[30]~93_combout ),
	.asdata(\_T_244[30]~53_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[30]~q ),
	.prn(vcc));
defparam \cycle[30] .is_wysiwyg = "true";
defparam \cycle[30] .power_up = "low";

cyclone10lp_lcell_comb \cycle[31]~95 (
	.dataa(\cycle[31]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\cycle[30]~94 ),
	.combout(\cycle[31]~95_combout ),
	.cout());
defparam \cycle[31]~95 .lut_mask = 16'h5A5A;
defparam \cycle[31]~95 .sum_lutc_input = "cin";

dffeas \cycle[31] (
	.clk(clock),
	.d(\cycle[31]~95_combout ),
	.asdata(\_T_246[31]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycle~36_combout ),
	.ena(vcc),
	.q(\cycle[31]~q ),
	.prn(vcc));
defparam \cycle[31] .is_wysiwyg = "true";
defparam \cycle[31] .power_up = "low";

cyclone10lp_lcell_comb \WideAnd1~0 (
	.dataa(\cycle[0]~q ),
	.datab(\cycle[1]~q ),
	.datac(\cycle[31]~q ),
	.datad(\cycle[30]~q ),
	.cin(gnd),
	.combout(\WideAnd1~0_combout ),
	.cout());
defparam \WideAnd1~0 .lut_mask = 16'h7FFF;
defparam \WideAnd1~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd1~1 (
	.dataa(\cycle[29]~q ),
	.datab(\cycle[28]~q ),
	.datac(\cycle[27]~q ),
	.datad(\cycle[26]~q ),
	.cin(gnd),
	.combout(\WideAnd1~1_combout ),
	.cout());
defparam \WideAnd1~1 .lut_mask = 16'h7FFF;
defparam \WideAnd1~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd1~2 (
	.dataa(\cycle[25]~q ),
	.datab(\cycle[24]~q ),
	.datac(\cycle[23]~q ),
	.datad(\cycle[22]~q ),
	.cin(gnd),
	.combout(\WideAnd1~2_combout ),
	.cout());
defparam \WideAnd1~2 .lut_mask = 16'h7FFF;
defparam \WideAnd1~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd1~3 (
	.dataa(\cycle[21]~q ),
	.datab(\cycle[20]~q ),
	.datac(\cycle[19]~q ),
	.datad(\cycle[18]~q ),
	.cin(gnd),
	.combout(\WideAnd1~3_combout ),
	.cout());
defparam \WideAnd1~3 .lut_mask = 16'h7FFF;
defparam \WideAnd1~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd1~4 (
	.dataa(\WideAnd1~0_combout ),
	.datab(\WideAnd1~1_combout ),
	.datac(\WideAnd1~2_combout ),
	.datad(\WideAnd1~3_combout ),
	.cin(gnd),
	.combout(\WideAnd1~4_combout ),
	.cout());
defparam \WideAnd1~4 .lut_mask = 16'hFFFE;
defparam \WideAnd1~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd1~5 (
	.dataa(\cycle[17]~q ),
	.datab(\cycle[16]~q ),
	.datac(\cycle[15]~q ),
	.datad(\cycle[14]~q ),
	.cin(gnd),
	.combout(\WideAnd1~5_combout ),
	.cout());
defparam \WideAnd1~5 .lut_mask = 16'h7FFF;
defparam \WideAnd1~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd1~6 (
	.dataa(\cycle[13]~q ),
	.datab(\cycle[12]~q ),
	.datac(\cycle[11]~q ),
	.datad(\cycle[10]~q ),
	.cin(gnd),
	.combout(\WideAnd1~6_combout ),
	.cout());
defparam \WideAnd1~6 .lut_mask = 16'h7FFF;
defparam \WideAnd1~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd1~7 (
	.dataa(\cycle[9]~q ),
	.datab(\cycle[8]~q ),
	.datac(\cycle[7]~q ),
	.datad(\cycle[6]~q ),
	.cin(gnd),
	.combout(\WideAnd1~7_combout ),
	.cout());
defparam \WideAnd1~7 .lut_mask = 16'h7FFF;
defparam \WideAnd1~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd1~8 (
	.dataa(\cycle[5]~q ),
	.datab(\cycle[4]~q ),
	.datac(\cycle[3]~q ),
	.datad(\cycle[2]~q ),
	.cin(gnd),
	.combout(\WideAnd1~8_combout ),
	.cout());
defparam \WideAnd1~8 .lut_mask = 16'h7FFF;
defparam \WideAnd1~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd1~9 (
	.dataa(\WideAnd1~5_combout ),
	.datab(\WideAnd1~6_combout ),
	.datac(\WideAnd1~7_combout ),
	.datad(\WideAnd1~8_combout ),
	.cin(gnd),
	.combout(\WideAnd1~9_combout ),
	.cout());
defparam \WideAnd1~9 .lut_mask = 16'hFFFE;
defparam \WideAnd1~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cycleh[23]~37 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\WideAnd1~4_combout ),
	.datac(\WideAnd1~9_combout ),
	.datad(\cycleh~36_combout ),
	.cin(gnd),
	.combout(\cycleh[23]~37_combout ),
	.cout());
defparam \cycleh[23]~37 .lut_mask = 16'hFF57;
defparam \cycleh[23]~37 .sum_lutc_input = "datac";

dffeas \cycleh[0] (
	.clk(clock),
	.d(\cycleh[0]~32_combout ),
	.asdata(\_T_246[0]~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[0]~q ),
	.prn(vcc));
defparam \cycleh[0] .is_wysiwyg = "true";
defparam \cycleh[0] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[1]~34 (
	.dataa(\cycleh[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[0]~33 ),
	.combout(\cycleh[1]~34_combout ),
	.cout(\cycleh[1]~35 ));
defparam \cycleh[1]~34 .lut_mask = 16'h5A5F;
defparam \cycleh[1]~34 .sum_lutc_input = "cin";

dffeas \cycleh[1] (
	.clk(clock),
	.d(\cycleh[1]~34_combout ),
	.asdata(\_T_246[1]~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[1]~q ),
	.prn(vcc));
defparam \cycleh[1] .is_wysiwyg = "true";
defparam \cycleh[1] .power_up = "low";

cyclone10lp_lcell_comb \mbadaddr[0]~0 (
	.dataa(\Equal28~0_combout ),
	.datab(\instreth~32_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mbadaddr[0]~0_combout ),
	.cout());
defparam \mbadaddr[0]~0 .lut_mask = 16'h8888;
defparam \mbadaddr[0]~0 .sum_lutc_input = "datac";

dffeas \mbadaddr[1] (
	.clk(clock),
	.d(\_T_246[1]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[1]~q ),
	.prn(vcc));
defparam \mbadaddr[1] .is_wysiwyg = "true";
defparam \mbadaddr[1] .power_up = "low";

cyclone10lp_lcell_comb \io_out[1]~11 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~10_combout ),
	.datac(\cycleh[1]~q ),
	.datad(\mbadaddr[1]~q ),
	.cin(gnd),
	.combout(\io_out[1]~11_combout ),
	.cout());
defparam \io_out[1]~11 .lut_mask = 16'hEAC0;
defparam \io_out[1]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \timeh~32 (
	.dataa(ex_csr_addr_6),
	.datab(\Equal23~0_combout ),
	.datac(ex_csr_addr_7),
	.datad(\Equal11~3_combout ),
	.cin(gnd),
	.combout(\timeh~32_combout ),
	.cout());
defparam \timeh~32 .lut_mask = 16'h0777;
defparam \timeh~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[1]~12 (
	.dataa(ex_csr_addr_7),
	.datab(\Equal4~0_combout ),
	.datac(\Equal3~0_combout ),
	.datad(\timeh~32_combout ),
	.cin(gnd),
	.combout(\io_out[1]~12_combout ),
	.cout());
defparam \io_out[1]~12 .lut_mask = 16'h80FF;
defparam \io_out[1]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \timeh[0]~34 (
	.dataa(\timeh[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\timeh[0]~34_combout ),
	.cout(\timeh[0]~35 ));
defparam \timeh[0]~34 .lut_mask = 16'h55AA;
defparam \timeh[0]~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \timeh~38 (
	.dataa(\timeh~33_combout ),
	.datab(ex_csr_addr_6),
	.datac(\Equal23~0_combout ),
	.datad(\timeh~32_combout ),
	.cin(gnd),
	.combout(\timeh~38_combout ),
	.cout());
defparam \timeh~38 .lut_mask = 16'h008A;
defparam \timeh~38 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \time_[2]~37 (
	.dataa(\time_[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[1]~35 ),
	.combout(\time_[2]~37_combout ),
	.cout(\time_[2]~38 ));
defparam \time_[2]~37 .lut_mask = 16'hA50A;
defparam \time_[2]~37 .sum_lutc_input = "cin";

dffeas \time_[2] (
	.clk(clock),
	.d(\time_[2]~37_combout ),
	.asdata(\_T_246[2]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[2]~q ),
	.prn(vcc));
defparam \time_[2] .is_wysiwyg = "true";
defparam \time_[2] .power_up = "low";

cyclone10lp_lcell_comb \time_[3]~39 (
	.dataa(\time_[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[2]~38 ),
	.combout(\time_[3]~39_combout ),
	.cout(\time_[3]~40 ));
defparam \time_[3]~39 .lut_mask = 16'h5A5F;
defparam \time_[3]~39 .sum_lutc_input = "cin";

dffeas \time_[3] (
	.clk(clock),
	.d(\time_[3]~39_combout ),
	.asdata(\_T_246[3]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[3]~q ),
	.prn(vcc));
defparam \time_[3] .is_wysiwyg = "true";
defparam \time_[3] .power_up = "low";

cyclone10lp_lcell_comb \time_[4]~41 (
	.dataa(\time_[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[3]~40 ),
	.combout(\time_[4]~41_combout ),
	.cout(\time_[4]~42 ));
defparam \time_[4]~41 .lut_mask = 16'hA50A;
defparam \time_[4]~41 .sum_lutc_input = "cin";

dffeas \time_[4] (
	.clk(clock),
	.d(\time_[4]~41_combout ),
	.asdata(\_T_244[4]~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[4]~q ),
	.prn(vcc));
defparam \time_[4] .is_wysiwyg = "true";
defparam \time_[4] .power_up = "low";

cyclone10lp_lcell_comb \time_[5]~43 (
	.dataa(\time_[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[4]~42 ),
	.combout(\time_[5]~43_combout ),
	.cout(\time_[5]~44 ));
defparam \time_[5]~43 .lut_mask = 16'h5A5F;
defparam \time_[5]~43 .sum_lutc_input = "cin";

dffeas \time_[5] (
	.clk(clock),
	.d(\time_[5]~43_combout ),
	.asdata(\_T_244[5]~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[5]~q ),
	.prn(vcc));
defparam \time_[5] .is_wysiwyg = "true";
defparam \time_[5] .power_up = "low";

cyclone10lp_lcell_comb \time_[6]~45 (
	.dataa(\time_[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[5]~44 ),
	.combout(\time_[6]~45_combout ),
	.cout(\time_[6]~46 ));
defparam \time_[6]~45 .lut_mask = 16'hA50A;
defparam \time_[6]~45 .sum_lutc_input = "cin";

dffeas \time_[6] (
	.clk(clock),
	.d(\time_[6]~45_combout ),
	.asdata(\_T_244[6]~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[6]~q ),
	.prn(vcc));
defparam \time_[6] .is_wysiwyg = "true";
defparam \time_[6] .power_up = "low";

cyclone10lp_lcell_comb \time_[7]~47 (
	.dataa(\time_[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[6]~46 ),
	.combout(\time_[7]~47_combout ),
	.cout(\time_[7]~48 ));
defparam \time_[7]~47 .lut_mask = 16'h5A5F;
defparam \time_[7]~47 .sum_lutc_input = "cin";

dffeas \time_[7] (
	.clk(clock),
	.d(\time_[7]~47_combout ),
	.asdata(\_T_244[7]~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[7]~q ),
	.prn(vcc));
defparam \time_[7] .is_wysiwyg = "true";
defparam \time_[7] .power_up = "low";

cyclone10lp_lcell_comb \time_[8]~49 (
	.dataa(\time_[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[7]~48 ),
	.combout(\time_[8]~49_combout ),
	.cout(\time_[8]~50 ));
defparam \time_[8]~49 .lut_mask = 16'hA50A;
defparam \time_[8]~49 .sum_lutc_input = "cin";

dffeas \time_[8] (
	.clk(clock),
	.d(\time_[8]~49_combout ),
	.asdata(\_T_244[8]~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[8]~q ),
	.prn(vcc));
defparam \time_[8] .is_wysiwyg = "true";
defparam \time_[8] .power_up = "low";

cyclone10lp_lcell_comb \time_[9]~51 (
	.dataa(\time_[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[8]~50 ),
	.combout(\time_[9]~51_combout ),
	.cout(\time_[9]~52 ));
defparam \time_[9]~51 .lut_mask = 16'h5A5F;
defparam \time_[9]~51 .sum_lutc_input = "cin";

dffeas \time_[9] (
	.clk(clock),
	.d(\time_[9]~51_combout ),
	.asdata(\_T_244[9]~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[9]~q ),
	.prn(vcc));
defparam \time_[9] .is_wysiwyg = "true";
defparam \time_[9] .power_up = "low";

cyclone10lp_lcell_comb \time_[10]~53 (
	.dataa(\time_[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[9]~52 ),
	.combout(\time_[10]~53_combout ),
	.cout(\time_[10]~54 ));
defparam \time_[10]~53 .lut_mask = 16'hA50A;
defparam \time_[10]~53 .sum_lutc_input = "cin";

dffeas \time_[10] (
	.clk(clock),
	.d(\time_[10]~53_combout ),
	.asdata(\_T_244[10]~13_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[10]~q ),
	.prn(vcc));
defparam \time_[10] .is_wysiwyg = "true";
defparam \time_[10] .power_up = "low";

cyclone10lp_lcell_comb \time_[11]~55 (
	.dataa(\time_[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[10]~54 ),
	.combout(\time_[11]~55_combout ),
	.cout(\time_[11]~56 ));
defparam \time_[11]~55 .lut_mask = 16'h5A5F;
defparam \time_[11]~55 .sum_lutc_input = "cin";

dffeas \time_[11] (
	.clk(clock),
	.d(\time_[11]~55_combout ),
	.asdata(\_T_244[11]~15_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[11]~q ),
	.prn(vcc));
defparam \time_[11] .is_wysiwyg = "true";
defparam \time_[11] .power_up = "low";

cyclone10lp_lcell_comb \time_[12]~57 (
	.dataa(\time_[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[11]~56 ),
	.combout(\time_[12]~57_combout ),
	.cout(\time_[12]~58 ));
defparam \time_[12]~57 .lut_mask = 16'hA50A;
defparam \time_[12]~57 .sum_lutc_input = "cin";

dffeas \time_[12] (
	.clk(clock),
	.d(\time_[12]~57_combout ),
	.asdata(\_T_244[12]~17_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[12]~q ),
	.prn(vcc));
defparam \time_[12] .is_wysiwyg = "true";
defparam \time_[12] .power_up = "low";

cyclone10lp_lcell_comb \time_[13]~59 (
	.dataa(\time_[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[12]~58 ),
	.combout(\time_[13]~59_combout ),
	.cout(\time_[13]~60 ));
defparam \time_[13]~59 .lut_mask = 16'h5A5F;
defparam \time_[13]~59 .sum_lutc_input = "cin";

dffeas \time_[13] (
	.clk(clock),
	.d(\time_[13]~59_combout ),
	.asdata(\_T_244[13]~19_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[13]~q ),
	.prn(vcc));
defparam \time_[13] .is_wysiwyg = "true";
defparam \time_[13] .power_up = "low";

cyclone10lp_lcell_comb \time_[14]~61 (
	.dataa(\time_[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[13]~60 ),
	.combout(\time_[14]~61_combout ),
	.cout(\time_[14]~62 ));
defparam \time_[14]~61 .lut_mask = 16'hA50A;
defparam \time_[14]~61 .sum_lutc_input = "cin";

dffeas \time_[14] (
	.clk(clock),
	.d(\time_[14]~61_combout ),
	.asdata(\_T_244[14]~21_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[14]~q ),
	.prn(vcc));
defparam \time_[14] .is_wysiwyg = "true";
defparam \time_[14] .power_up = "low";

cyclone10lp_lcell_comb \time_[15]~63 (
	.dataa(\time_[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[14]~62 ),
	.combout(\time_[15]~63_combout ),
	.cout(\time_[15]~64 ));
defparam \time_[15]~63 .lut_mask = 16'h5A5F;
defparam \time_[15]~63 .sum_lutc_input = "cin";

dffeas \time_[15] (
	.clk(clock),
	.d(\time_[15]~63_combout ),
	.asdata(\_T_244[15]~23_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[15]~q ),
	.prn(vcc));
defparam \time_[15] .is_wysiwyg = "true";
defparam \time_[15] .power_up = "low";

cyclone10lp_lcell_comb \time_[16]~65 (
	.dataa(\time_[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[15]~64 ),
	.combout(\time_[16]~65_combout ),
	.cout(\time_[16]~66 ));
defparam \time_[16]~65 .lut_mask = 16'hA50A;
defparam \time_[16]~65 .sum_lutc_input = "cin";

dffeas \time_[16] (
	.clk(clock),
	.d(\time_[16]~65_combout ),
	.asdata(\_T_244[16]~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[16]~q ),
	.prn(vcc));
defparam \time_[16] .is_wysiwyg = "true";
defparam \time_[16] .power_up = "low";

cyclone10lp_lcell_comb \time_[17]~67 (
	.dataa(\time_[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[16]~66 ),
	.combout(\time_[17]~67_combout ),
	.cout(\time_[17]~68 ));
defparam \time_[17]~67 .lut_mask = 16'h5A5F;
defparam \time_[17]~67 .sum_lutc_input = "cin";

dffeas \time_[17] (
	.clk(clock),
	.d(\time_[17]~67_combout ),
	.asdata(\_T_244[17]~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[17]~q ),
	.prn(vcc));
defparam \time_[17] .is_wysiwyg = "true";
defparam \time_[17] .power_up = "low";

cyclone10lp_lcell_comb \time_[18]~69 (
	.dataa(\time_[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[17]~68 ),
	.combout(\time_[18]~69_combout ),
	.cout(\time_[18]~70 ));
defparam \time_[18]~69 .lut_mask = 16'hA50A;
defparam \time_[18]~69 .sum_lutc_input = "cin";

dffeas \time_[18] (
	.clk(clock),
	.d(\time_[18]~69_combout ),
	.asdata(\_T_244[18]~29_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[18]~q ),
	.prn(vcc));
defparam \time_[18] .is_wysiwyg = "true";
defparam \time_[18] .power_up = "low";

cyclone10lp_lcell_comb \time_[19]~71 (
	.dataa(\time_[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[18]~70 ),
	.combout(\time_[19]~71_combout ),
	.cout(\time_[19]~72 ));
defparam \time_[19]~71 .lut_mask = 16'h5A5F;
defparam \time_[19]~71 .sum_lutc_input = "cin";

dffeas \time_[19] (
	.clk(clock),
	.d(\time_[19]~71_combout ),
	.asdata(\_T_244[19]~31_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[19]~q ),
	.prn(vcc));
defparam \time_[19] .is_wysiwyg = "true";
defparam \time_[19] .power_up = "low";

cyclone10lp_lcell_comb \time_[20]~73 (
	.dataa(\time_[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[19]~72 ),
	.combout(\time_[20]~73_combout ),
	.cout(\time_[20]~74 ));
defparam \time_[20]~73 .lut_mask = 16'hA50A;
defparam \time_[20]~73 .sum_lutc_input = "cin";

dffeas \time_[20] (
	.clk(clock),
	.d(\time_[20]~73_combout ),
	.asdata(\_T_244[20]~33_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[20]~q ),
	.prn(vcc));
defparam \time_[20] .is_wysiwyg = "true";
defparam \time_[20] .power_up = "low";

cyclone10lp_lcell_comb \time_[21]~75 (
	.dataa(\time_[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[20]~74 ),
	.combout(\time_[21]~75_combout ),
	.cout(\time_[21]~76 ));
defparam \time_[21]~75 .lut_mask = 16'h5A5F;
defparam \time_[21]~75 .sum_lutc_input = "cin";

dffeas \time_[21] (
	.clk(clock),
	.d(\time_[21]~75_combout ),
	.asdata(\_T_244[21]~35_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[21]~q ),
	.prn(vcc));
defparam \time_[21] .is_wysiwyg = "true";
defparam \time_[21] .power_up = "low";

cyclone10lp_lcell_comb \time_[22]~77 (
	.dataa(\time_[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[21]~76 ),
	.combout(\time_[22]~77_combout ),
	.cout(\time_[22]~78 ));
defparam \time_[22]~77 .lut_mask = 16'hA50A;
defparam \time_[22]~77 .sum_lutc_input = "cin";

dffeas \time_[22] (
	.clk(clock),
	.d(\time_[22]~77_combout ),
	.asdata(\_T_244[22]~37_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[22]~q ),
	.prn(vcc));
defparam \time_[22] .is_wysiwyg = "true";
defparam \time_[22] .power_up = "low";

cyclone10lp_lcell_comb \time_[23]~79 (
	.dataa(\time_[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[22]~78 ),
	.combout(\time_[23]~79_combout ),
	.cout(\time_[23]~80 ));
defparam \time_[23]~79 .lut_mask = 16'h5A5F;
defparam \time_[23]~79 .sum_lutc_input = "cin";

dffeas \time_[23] (
	.clk(clock),
	.d(\time_[23]~79_combout ),
	.asdata(\_T_244[23]~39_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[23]~q ),
	.prn(vcc));
defparam \time_[23] .is_wysiwyg = "true";
defparam \time_[23] .power_up = "low";

cyclone10lp_lcell_comb \time_[24]~81 (
	.dataa(\time_[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[23]~80 ),
	.combout(\time_[24]~81_combout ),
	.cout(\time_[24]~82 ));
defparam \time_[24]~81 .lut_mask = 16'hA50A;
defparam \time_[24]~81 .sum_lutc_input = "cin";

dffeas \time_[24] (
	.clk(clock),
	.d(\time_[24]~81_combout ),
	.asdata(\_T_244[24]~41_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[24]~q ),
	.prn(vcc));
defparam \time_[24] .is_wysiwyg = "true";
defparam \time_[24] .power_up = "low";

cyclone10lp_lcell_comb \time_[25]~83 (
	.dataa(\time_[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[24]~82 ),
	.combout(\time_[25]~83_combout ),
	.cout(\time_[25]~84 ));
defparam \time_[25]~83 .lut_mask = 16'h5A5F;
defparam \time_[25]~83 .sum_lutc_input = "cin";

dffeas \time_[25] (
	.clk(clock),
	.d(\time_[25]~83_combout ),
	.asdata(\_T_244[25]~43_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[25]~q ),
	.prn(vcc));
defparam \time_[25] .is_wysiwyg = "true";
defparam \time_[25] .power_up = "low";

cyclone10lp_lcell_comb \time_[26]~85 (
	.dataa(\time_[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[25]~84 ),
	.combout(\time_[26]~85_combout ),
	.cout(\time_[26]~86 ));
defparam \time_[26]~85 .lut_mask = 16'hA50A;
defparam \time_[26]~85 .sum_lutc_input = "cin";

dffeas \time_[26] (
	.clk(clock),
	.d(\time_[26]~85_combout ),
	.asdata(\_T_244[26]~45_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[26]~q ),
	.prn(vcc));
defparam \time_[26] .is_wysiwyg = "true";
defparam \time_[26] .power_up = "low";

cyclone10lp_lcell_comb \time_[27]~87 (
	.dataa(\time_[27]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[26]~86 ),
	.combout(\time_[27]~87_combout ),
	.cout(\time_[27]~88 ));
defparam \time_[27]~87 .lut_mask = 16'h5A5F;
defparam \time_[27]~87 .sum_lutc_input = "cin";

dffeas \time_[27] (
	.clk(clock),
	.d(\time_[27]~87_combout ),
	.asdata(\_T_244[27]~47_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[27]~q ),
	.prn(vcc));
defparam \time_[27] .is_wysiwyg = "true";
defparam \time_[27] .power_up = "low";

cyclone10lp_lcell_comb \time_[28]~89 (
	.dataa(\time_[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[27]~88 ),
	.combout(\time_[28]~89_combout ),
	.cout(\time_[28]~90 ));
defparam \time_[28]~89 .lut_mask = 16'hA50A;
defparam \time_[28]~89 .sum_lutc_input = "cin";

dffeas \time_[28] (
	.clk(clock),
	.d(\time_[28]~89_combout ),
	.asdata(\_T_244[28]~49_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[28]~q ),
	.prn(vcc));
defparam \time_[28] .is_wysiwyg = "true";
defparam \time_[28] .power_up = "low";

cyclone10lp_lcell_comb \time_[29]~91 (
	.dataa(\time_[29]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[28]~90 ),
	.combout(\time_[29]~91_combout ),
	.cout(\time_[29]~92 ));
defparam \time_[29]~91 .lut_mask = 16'h5A5F;
defparam \time_[29]~91 .sum_lutc_input = "cin";

dffeas \time_[29] (
	.clk(clock),
	.d(\time_[29]~91_combout ),
	.asdata(\_T_244[29]~51_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[29]~q ),
	.prn(vcc));
defparam \time_[29] .is_wysiwyg = "true";
defparam \time_[29] .power_up = "low";

cyclone10lp_lcell_comb \time_[30]~93 (
	.dataa(\time_[30]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\time_[29]~92 ),
	.combout(\time_[30]~93_combout ),
	.cout(\time_[30]~94 ));
defparam \time_[30]~93 .lut_mask = 16'hA50A;
defparam \time_[30]~93 .sum_lutc_input = "cin";

dffeas \time_[30] (
	.clk(clock),
	.d(\time_[30]~93_combout ),
	.asdata(\_T_244[30]~53_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[30]~q ),
	.prn(vcc));
defparam \time_[30] .is_wysiwyg = "true";
defparam \time_[30] .power_up = "low";

cyclone10lp_lcell_comb \time_[31]~95 (
	.dataa(\time_[31]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\time_[30]~94 ),
	.combout(\time_[31]~95_combout ),
	.cout());
defparam \time_[31]~95 .lut_mask = 16'h5A5A;
defparam \time_[31]~95 .sum_lutc_input = "cin";

dffeas \time_[31] (
	.clk(clock),
	.d(\time_[31]~95_combout ),
	.asdata(\_T_246[31]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\time_~36_combout ),
	.ena(vcc),
	.q(\time_[31]~q ),
	.prn(vcc));
defparam \time_[31] .is_wysiwyg = "true";
defparam \time_[31] .power_up = "low";

cyclone10lp_lcell_comb \WideAnd0~0 (
	.dataa(\time_[0]~q ),
	.datab(\time_[1]~q ),
	.datac(\time_[31]~q ),
	.datad(\time_[30]~q ),
	.cin(gnd),
	.combout(\WideAnd0~0_combout ),
	.cout());
defparam \WideAnd0~0 .lut_mask = 16'h7FFF;
defparam \WideAnd0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd0~1 (
	.dataa(\time_[29]~q ),
	.datab(\time_[28]~q ),
	.datac(\time_[27]~q ),
	.datad(\time_[26]~q ),
	.cin(gnd),
	.combout(\WideAnd0~1_combout ),
	.cout());
defparam \WideAnd0~1 .lut_mask = 16'h7FFF;
defparam \WideAnd0~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd0~2 (
	.dataa(\time_[25]~q ),
	.datab(\time_[24]~q ),
	.datac(\time_[23]~q ),
	.datad(\time_[22]~q ),
	.cin(gnd),
	.combout(\WideAnd0~2_combout ),
	.cout());
defparam \WideAnd0~2 .lut_mask = 16'h7FFF;
defparam \WideAnd0~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd0~3 (
	.dataa(\time_[21]~q ),
	.datab(\time_[20]~q ),
	.datac(\time_[19]~q ),
	.datad(\time_[18]~q ),
	.cin(gnd),
	.combout(\WideAnd0~3_combout ),
	.cout());
defparam \WideAnd0~3 .lut_mask = 16'h7FFF;
defparam \WideAnd0~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd0~4 (
	.dataa(\WideAnd0~0_combout ),
	.datab(\WideAnd0~1_combout ),
	.datac(\WideAnd0~2_combout ),
	.datad(\WideAnd0~3_combout ),
	.cin(gnd),
	.combout(\WideAnd0~4_combout ),
	.cout());
defparam \WideAnd0~4 .lut_mask = 16'hFFFE;
defparam \WideAnd0~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd0~5 (
	.dataa(\time_[17]~q ),
	.datab(\time_[16]~q ),
	.datac(\time_[15]~q ),
	.datad(\time_[14]~q ),
	.cin(gnd),
	.combout(\WideAnd0~5_combout ),
	.cout());
defparam \WideAnd0~5 .lut_mask = 16'h7FFF;
defparam \WideAnd0~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd0~6 (
	.dataa(\time_[13]~q ),
	.datab(\time_[12]~q ),
	.datac(\time_[11]~q ),
	.datad(\time_[10]~q ),
	.cin(gnd),
	.combout(\WideAnd0~6_combout ),
	.cout());
defparam \WideAnd0~6 .lut_mask = 16'h7FFF;
defparam \WideAnd0~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd0~7 (
	.dataa(\time_[9]~q ),
	.datab(\time_[8]~q ),
	.datac(\time_[7]~q ),
	.datad(\time_[6]~q ),
	.cin(gnd),
	.combout(\WideAnd0~7_combout ),
	.cout());
defparam \WideAnd0~7 .lut_mask = 16'h7FFF;
defparam \WideAnd0~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd0~8 (
	.dataa(\time_[5]~q ),
	.datab(\time_[4]~q ),
	.datac(\time_[3]~q ),
	.datad(\time_[2]~q ),
	.cin(gnd),
	.combout(\WideAnd0~8_combout ),
	.cout());
defparam \WideAnd0~8 .lut_mask = 16'h7FFF;
defparam \WideAnd0~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \WideAnd0~9 (
	.dataa(\WideAnd0~5_combout ),
	.datab(\WideAnd0~6_combout ),
	.datac(\WideAnd0~7_combout ),
	.datad(\WideAnd0~8_combout ),
	.cin(gnd),
	.combout(\WideAnd0~9_combout ),
	.cout());
defparam \WideAnd0~9 .lut_mask = 16'hFFFE;
defparam \WideAnd0~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \timeh[31]~39 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\WideAnd0~4_combout ),
	.datac(\WideAnd0~9_combout ),
	.datad(\timeh~38_combout ),
	.cin(gnd),
	.combout(\timeh[31]~39_combout ),
	.cout());
defparam \timeh[31]~39 .lut_mask = 16'hFF57;
defparam \timeh[31]~39 .sum_lutc_input = "datac";

dffeas \timeh[0] (
	.clk(clock),
	.d(\timeh[0]~34_combout ),
	.asdata(\_T_246[0]~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[0]~q ),
	.prn(vcc));
defparam \timeh[0] .is_wysiwyg = "true";
defparam \timeh[0] .power_up = "low";

cyclone10lp_lcell_comb \timeh[1]~36 (
	.dataa(\timeh[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[0]~35 ),
	.combout(\timeh[1]~36_combout ),
	.cout(\timeh[1]~37 ));
defparam \timeh[1]~36 .lut_mask = 16'h5A5F;
defparam \timeh[1]~36 .sum_lutc_input = "cin";

dffeas \timeh[1] (
	.clk(clock),
	.d(\timeh[1]~36_combout ),
	.asdata(\_T_246[1]~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[1]~q ),
	.prn(vcc));
defparam \timeh[1] .is_wysiwyg = "true";
defparam \timeh[1] .power_up = "low";

cyclone10lp_lcell_comb \io_out[1]~13 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_1),
	.datad(\timeh[1]~q ),
	.cin(gnd),
	.combout(\io_out[1]~13_combout ),
	.cout());
defparam \io_out[1]~13 .lut_mask = 16'hEAC0;
defparam \io_out[1]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal13~1 (
	.dataa(ex_csr_addr_7),
	.datab(\Equal11~2_combout ),
	.datac(gnd),
	.datad(ex_csr_addr_0),
	.cin(gnd),
	.combout(\Equal13~1_combout ),
	.cout());
defparam \Equal13~1 .lut_mask = 16'h0088;
defparam \Equal13~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[1]~14 (
	.dataa(ex_csr_addr_1),
	.datab(ex_csr_addr_7),
	.datac(\Equal8~0_combout ),
	.datad(\Equal13~1_combout ),
	.cin(gnd),
	.combout(\io_out[1]~14_combout ),
	.cout());
defparam \io_out[1]~14 .lut_mask = 16'hEAC0;
defparam \io_out[1]~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \instreth[0]~33 (
	.dataa(\instreth[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\instreth[0]~33_combout ),
	.cout(\instreth[0]~34 ));
defparam \instreth[0]~33 .lut_mask = 16'h55AA;
defparam \instreth[0]~33 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \instreth~37 (
	.dataa(\Equal13~1_combout ),
	.datab(\instreth~32_combout ),
	.datac(gnd),
	.datad(\Equal13~0_combout ),
	.cin(gnd),
	.combout(\instreth~37_combout ),
	.cout());
defparam \instreth~37 .lut_mask = 16'h0088;
defparam \instreth~37 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb isInstRet(
	.dataa(\isInstRet~0_combout ),
	.datab(gnd),
	.datac(io_expt1),
	.datad(isEcall),
	.cin(gnd),
	.combout(\isInstRet~combout ),
	.cout());
defparam isInstRet.lut_mask = 16'hAAAF;
defparam isInstRet.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \instret[2]~39 (
	.dataa(\instret[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[1]~37 ),
	.combout(\instret[2]~39_combout ),
	.cout(\instret[2]~40 ));
defparam \instret[2]~39 .lut_mask = 16'hA50A;
defparam \instret[2]~39 .sum_lutc_input = "cin";

dffeas \instret[2] (
	.clk(clock),
	.d(\instret[2]~39_combout ),
	.asdata(\_T_246[2]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[2]~q ),
	.prn(vcc));
defparam \instret[2] .is_wysiwyg = "true";
defparam \instret[2] .power_up = "low";

cyclone10lp_lcell_comb \instret[3]~41 (
	.dataa(\instret[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[2]~40 ),
	.combout(\instret[3]~41_combout ),
	.cout(\instret[3]~42 ));
defparam \instret[3]~41 .lut_mask = 16'h5A5F;
defparam \instret[3]~41 .sum_lutc_input = "cin";

dffeas \instret[3] (
	.clk(clock),
	.d(\instret[3]~41_combout ),
	.asdata(\_T_246[3]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[3]~q ),
	.prn(vcc));
defparam \instret[3] .is_wysiwyg = "true";
defparam \instret[3] .power_up = "low";

cyclone10lp_lcell_comb \instret[4]~43 (
	.dataa(\instret[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[3]~42 ),
	.combout(\instret[4]~43_combout ),
	.cout(\instret[4]~44 ));
defparam \instret[4]~43 .lut_mask = 16'hA50A;
defparam \instret[4]~43 .sum_lutc_input = "cin";

dffeas \instret[4] (
	.clk(clock),
	.d(\instret[4]~43_combout ),
	.asdata(\_T_244[4]~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[4]~q ),
	.prn(vcc));
defparam \instret[4] .is_wysiwyg = "true";
defparam \instret[4] .power_up = "low";

cyclone10lp_lcell_comb \instret[5]~45 (
	.dataa(\instret[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[4]~44 ),
	.combout(\instret[5]~45_combout ),
	.cout(\instret[5]~46 ));
defparam \instret[5]~45 .lut_mask = 16'h5A5F;
defparam \instret[5]~45 .sum_lutc_input = "cin";

dffeas \instret[5] (
	.clk(clock),
	.d(\instret[5]~45_combout ),
	.asdata(\_T_244[5]~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[5]~q ),
	.prn(vcc));
defparam \instret[5] .is_wysiwyg = "true";
defparam \instret[5] .power_up = "low";

cyclone10lp_lcell_comb \instret[6]~47 (
	.dataa(\instret[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[5]~46 ),
	.combout(\instret[6]~47_combout ),
	.cout(\instret[6]~48 ));
defparam \instret[6]~47 .lut_mask = 16'hA50A;
defparam \instret[6]~47 .sum_lutc_input = "cin";

dffeas \instret[6] (
	.clk(clock),
	.d(\instret[6]~47_combout ),
	.asdata(\_T_244[6]~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[6]~q ),
	.prn(vcc));
defparam \instret[6] .is_wysiwyg = "true";
defparam \instret[6] .power_up = "low";

cyclone10lp_lcell_comb \instret[7]~49 (
	.dataa(\instret[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[6]~48 ),
	.combout(\instret[7]~49_combout ),
	.cout(\instret[7]~50 ));
defparam \instret[7]~49 .lut_mask = 16'h5A5F;
defparam \instret[7]~49 .sum_lutc_input = "cin";

dffeas \instret[7] (
	.clk(clock),
	.d(\instret[7]~49_combout ),
	.asdata(\_T_244[7]~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[7]~q ),
	.prn(vcc));
defparam \instret[7] .is_wysiwyg = "true";
defparam \instret[7] .power_up = "low";

cyclone10lp_lcell_comb \instret[8]~51 (
	.dataa(\instret[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[7]~50 ),
	.combout(\instret[8]~51_combout ),
	.cout(\instret[8]~52 ));
defparam \instret[8]~51 .lut_mask = 16'hA50A;
defparam \instret[8]~51 .sum_lutc_input = "cin";

dffeas \instret[8] (
	.clk(clock),
	.d(\instret[8]~51_combout ),
	.asdata(\_T_244[8]~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[8]~q ),
	.prn(vcc));
defparam \instret[8] .is_wysiwyg = "true";
defparam \instret[8] .power_up = "low";

cyclone10lp_lcell_comb \instret[9]~53 (
	.dataa(\instret[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[8]~52 ),
	.combout(\instret[9]~53_combout ),
	.cout(\instret[9]~54 ));
defparam \instret[9]~53 .lut_mask = 16'h5A5F;
defparam \instret[9]~53 .sum_lutc_input = "cin";

dffeas \instret[9] (
	.clk(clock),
	.d(\instret[9]~53_combout ),
	.asdata(\_T_244[9]~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[9]~q ),
	.prn(vcc));
defparam \instret[9] .is_wysiwyg = "true";
defparam \instret[9] .power_up = "low";

cyclone10lp_lcell_comb \instret[10]~55 (
	.dataa(\instret[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[9]~54 ),
	.combout(\instret[10]~55_combout ),
	.cout(\instret[10]~56 ));
defparam \instret[10]~55 .lut_mask = 16'hA50A;
defparam \instret[10]~55 .sum_lutc_input = "cin";

dffeas \instret[10] (
	.clk(clock),
	.d(\instret[10]~55_combout ),
	.asdata(\_T_244[10]~13_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[10]~q ),
	.prn(vcc));
defparam \instret[10] .is_wysiwyg = "true";
defparam \instret[10] .power_up = "low";

cyclone10lp_lcell_comb \instret[11]~57 (
	.dataa(\instret[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[10]~56 ),
	.combout(\instret[11]~57_combout ),
	.cout(\instret[11]~58 ));
defparam \instret[11]~57 .lut_mask = 16'h5A5F;
defparam \instret[11]~57 .sum_lutc_input = "cin";

dffeas \instret[11] (
	.clk(clock),
	.d(\instret[11]~57_combout ),
	.asdata(\_T_244[11]~15_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[11]~q ),
	.prn(vcc));
defparam \instret[11] .is_wysiwyg = "true";
defparam \instret[11] .power_up = "low";

cyclone10lp_lcell_comb \instret[12]~59 (
	.dataa(\instret[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[11]~58 ),
	.combout(\instret[12]~59_combout ),
	.cout(\instret[12]~60 ));
defparam \instret[12]~59 .lut_mask = 16'hA50A;
defparam \instret[12]~59 .sum_lutc_input = "cin";

dffeas \instret[12] (
	.clk(clock),
	.d(\instret[12]~59_combout ),
	.asdata(\_T_244[12]~17_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[12]~q ),
	.prn(vcc));
defparam \instret[12] .is_wysiwyg = "true";
defparam \instret[12] .power_up = "low";

cyclone10lp_lcell_comb \instret[13]~61 (
	.dataa(\instret[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[12]~60 ),
	.combout(\instret[13]~61_combout ),
	.cout(\instret[13]~62 ));
defparam \instret[13]~61 .lut_mask = 16'h5A5F;
defparam \instret[13]~61 .sum_lutc_input = "cin";

dffeas \instret[13] (
	.clk(clock),
	.d(\instret[13]~61_combout ),
	.asdata(\_T_244[13]~19_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[13]~q ),
	.prn(vcc));
defparam \instret[13] .is_wysiwyg = "true";
defparam \instret[13] .power_up = "low";

cyclone10lp_lcell_comb \instret[14]~63 (
	.dataa(\instret[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[13]~62 ),
	.combout(\instret[14]~63_combout ),
	.cout(\instret[14]~64 ));
defparam \instret[14]~63 .lut_mask = 16'hA50A;
defparam \instret[14]~63 .sum_lutc_input = "cin";

dffeas \instret[14] (
	.clk(clock),
	.d(\instret[14]~63_combout ),
	.asdata(\_T_244[14]~21_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[14]~q ),
	.prn(vcc));
defparam \instret[14] .is_wysiwyg = "true";
defparam \instret[14] .power_up = "low";

cyclone10lp_lcell_comb \instret[15]~65 (
	.dataa(\instret[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[14]~64 ),
	.combout(\instret[15]~65_combout ),
	.cout(\instret[15]~66 ));
defparam \instret[15]~65 .lut_mask = 16'h5A5F;
defparam \instret[15]~65 .sum_lutc_input = "cin";

dffeas \instret[15] (
	.clk(clock),
	.d(\instret[15]~65_combout ),
	.asdata(\_T_244[15]~23_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[15]~q ),
	.prn(vcc));
defparam \instret[15] .is_wysiwyg = "true";
defparam \instret[15] .power_up = "low";

cyclone10lp_lcell_comb \instret[16]~67 (
	.dataa(\instret[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[15]~66 ),
	.combout(\instret[16]~67_combout ),
	.cout(\instret[16]~68 ));
defparam \instret[16]~67 .lut_mask = 16'hA50A;
defparam \instret[16]~67 .sum_lutc_input = "cin";

dffeas \instret[16] (
	.clk(clock),
	.d(\instret[16]~67_combout ),
	.asdata(\_T_244[16]~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[16]~q ),
	.prn(vcc));
defparam \instret[16] .is_wysiwyg = "true";
defparam \instret[16] .power_up = "low";

cyclone10lp_lcell_comb \instret[17]~69 (
	.dataa(\instret[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[16]~68 ),
	.combout(\instret[17]~69_combout ),
	.cout(\instret[17]~70 ));
defparam \instret[17]~69 .lut_mask = 16'h5A5F;
defparam \instret[17]~69 .sum_lutc_input = "cin";

dffeas \instret[17] (
	.clk(clock),
	.d(\instret[17]~69_combout ),
	.asdata(\_T_244[17]~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[17]~q ),
	.prn(vcc));
defparam \instret[17] .is_wysiwyg = "true";
defparam \instret[17] .power_up = "low";

cyclone10lp_lcell_comb \instret[18]~71 (
	.dataa(\instret[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[17]~70 ),
	.combout(\instret[18]~71_combout ),
	.cout(\instret[18]~72 ));
defparam \instret[18]~71 .lut_mask = 16'hA50A;
defparam \instret[18]~71 .sum_lutc_input = "cin";

dffeas \instret[18] (
	.clk(clock),
	.d(\instret[18]~71_combout ),
	.asdata(\_T_244[18]~29_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[18]~q ),
	.prn(vcc));
defparam \instret[18] .is_wysiwyg = "true";
defparam \instret[18] .power_up = "low";

cyclone10lp_lcell_comb \instret[19]~73 (
	.dataa(\instret[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[18]~72 ),
	.combout(\instret[19]~73_combout ),
	.cout(\instret[19]~74 ));
defparam \instret[19]~73 .lut_mask = 16'h5A5F;
defparam \instret[19]~73 .sum_lutc_input = "cin";

dffeas \instret[19] (
	.clk(clock),
	.d(\instret[19]~73_combout ),
	.asdata(\_T_244[19]~31_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[19]~q ),
	.prn(vcc));
defparam \instret[19] .is_wysiwyg = "true";
defparam \instret[19] .power_up = "low";

cyclone10lp_lcell_comb \instret[20]~75 (
	.dataa(\instret[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[19]~74 ),
	.combout(\instret[20]~75_combout ),
	.cout(\instret[20]~76 ));
defparam \instret[20]~75 .lut_mask = 16'hA50A;
defparam \instret[20]~75 .sum_lutc_input = "cin";

dffeas \instret[20] (
	.clk(clock),
	.d(\instret[20]~75_combout ),
	.asdata(\_T_244[20]~33_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[20]~q ),
	.prn(vcc));
defparam \instret[20] .is_wysiwyg = "true";
defparam \instret[20] .power_up = "low";

cyclone10lp_lcell_comb \instret[21]~77 (
	.dataa(\instret[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[20]~76 ),
	.combout(\instret[21]~77_combout ),
	.cout(\instret[21]~78 ));
defparam \instret[21]~77 .lut_mask = 16'h5A5F;
defparam \instret[21]~77 .sum_lutc_input = "cin";

dffeas \instret[21] (
	.clk(clock),
	.d(\instret[21]~77_combout ),
	.asdata(\_T_244[21]~35_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[21]~q ),
	.prn(vcc));
defparam \instret[21] .is_wysiwyg = "true";
defparam \instret[21] .power_up = "low";

cyclone10lp_lcell_comb \instret[22]~79 (
	.dataa(\instret[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[21]~78 ),
	.combout(\instret[22]~79_combout ),
	.cout(\instret[22]~80 ));
defparam \instret[22]~79 .lut_mask = 16'hA50A;
defparam \instret[22]~79 .sum_lutc_input = "cin";

dffeas \instret[22] (
	.clk(clock),
	.d(\instret[22]~79_combout ),
	.asdata(\_T_244[22]~37_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[22]~q ),
	.prn(vcc));
defparam \instret[22] .is_wysiwyg = "true";
defparam \instret[22] .power_up = "low";

cyclone10lp_lcell_comb \instret[23]~81 (
	.dataa(\instret[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[22]~80 ),
	.combout(\instret[23]~81_combout ),
	.cout(\instret[23]~82 ));
defparam \instret[23]~81 .lut_mask = 16'h5A5F;
defparam \instret[23]~81 .sum_lutc_input = "cin";

dffeas \instret[23] (
	.clk(clock),
	.d(\instret[23]~81_combout ),
	.asdata(\_T_244[23]~39_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[23]~q ),
	.prn(vcc));
defparam \instret[23] .is_wysiwyg = "true";
defparam \instret[23] .power_up = "low";

cyclone10lp_lcell_comb \instret[24]~83 (
	.dataa(\instret[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[23]~82 ),
	.combout(\instret[24]~83_combout ),
	.cout(\instret[24]~84 ));
defparam \instret[24]~83 .lut_mask = 16'hA50A;
defparam \instret[24]~83 .sum_lutc_input = "cin";

dffeas \instret[24] (
	.clk(clock),
	.d(\instret[24]~83_combout ),
	.asdata(\_T_244[24]~41_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[24]~q ),
	.prn(vcc));
defparam \instret[24] .is_wysiwyg = "true";
defparam \instret[24] .power_up = "low";

cyclone10lp_lcell_comb \instret[25]~85 (
	.dataa(\instret[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[24]~84 ),
	.combout(\instret[25]~85_combout ),
	.cout(\instret[25]~86 ));
defparam \instret[25]~85 .lut_mask = 16'h5A5F;
defparam \instret[25]~85 .sum_lutc_input = "cin";

dffeas \instret[25] (
	.clk(clock),
	.d(\instret[25]~85_combout ),
	.asdata(\_T_244[25]~43_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[25]~q ),
	.prn(vcc));
defparam \instret[25] .is_wysiwyg = "true";
defparam \instret[25] .power_up = "low";

cyclone10lp_lcell_comb \instret[26]~87 (
	.dataa(\instret[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[25]~86 ),
	.combout(\instret[26]~87_combout ),
	.cout(\instret[26]~88 ));
defparam \instret[26]~87 .lut_mask = 16'hA50A;
defparam \instret[26]~87 .sum_lutc_input = "cin";

dffeas \instret[26] (
	.clk(clock),
	.d(\instret[26]~87_combout ),
	.asdata(\_T_244[26]~45_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[26]~q ),
	.prn(vcc));
defparam \instret[26] .is_wysiwyg = "true";
defparam \instret[26] .power_up = "low";

cyclone10lp_lcell_comb \instret[27]~89 (
	.dataa(\instret[27]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[26]~88 ),
	.combout(\instret[27]~89_combout ),
	.cout(\instret[27]~90 ));
defparam \instret[27]~89 .lut_mask = 16'h5A5F;
defparam \instret[27]~89 .sum_lutc_input = "cin";

dffeas \instret[27] (
	.clk(clock),
	.d(\instret[27]~89_combout ),
	.asdata(\_T_244[27]~47_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[27]~q ),
	.prn(vcc));
defparam \instret[27] .is_wysiwyg = "true";
defparam \instret[27] .power_up = "low";

cyclone10lp_lcell_comb \instret[28]~91 (
	.dataa(\instret[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[27]~90 ),
	.combout(\instret[28]~91_combout ),
	.cout(\instret[28]~92 ));
defparam \instret[28]~91 .lut_mask = 16'hA50A;
defparam \instret[28]~91 .sum_lutc_input = "cin";

dffeas \instret[28] (
	.clk(clock),
	.d(\instret[28]~91_combout ),
	.asdata(\_T_244[28]~49_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[28]~q ),
	.prn(vcc));
defparam \instret[28] .is_wysiwyg = "true";
defparam \instret[28] .power_up = "low";

cyclone10lp_lcell_comb \instret[29]~93 (
	.dataa(\instret[29]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[28]~92 ),
	.combout(\instret[29]~93_combout ),
	.cout(\instret[29]~94 ));
defparam \instret[29]~93 .lut_mask = 16'h5A5F;
defparam \instret[29]~93 .sum_lutc_input = "cin";

dffeas \instret[29] (
	.clk(clock),
	.d(\instret[29]~93_combout ),
	.asdata(\_T_244[29]~51_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[29]~q ),
	.prn(vcc));
defparam \instret[29] .is_wysiwyg = "true";
defparam \instret[29] .power_up = "low";

cyclone10lp_lcell_comb \instret[30]~95 (
	.dataa(\instret[30]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instret[29]~94 ),
	.combout(\instret[30]~95_combout ),
	.cout(\instret[30]~96 ));
defparam \instret[30]~95 .lut_mask = 16'hA50A;
defparam \instret[30]~95 .sum_lutc_input = "cin";

dffeas \instret[30] (
	.clk(clock),
	.d(\instret[30]~95_combout ),
	.asdata(\_T_244[30]~53_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[30]~q ),
	.prn(vcc));
defparam \instret[30] .is_wysiwyg = "true";
defparam \instret[30] .power_up = "low";

cyclone10lp_lcell_comb \instret[31]~97 (
	.dataa(\instret[31]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\instret[30]~96 ),
	.combout(\instret[31]~97_combout ),
	.cout());
defparam \instret[31]~97 .lut_mask = 16'h5A5A;
defparam \instret[31]~97 .sum_lutc_input = "cin";

dffeas \instret[31] (
	.clk(clock),
	.d(\instret[31]~97_combout ),
	.asdata(\_T_246[31]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instret~38_combout ),
	.ena(\instret[0]~99_combout ),
	.q(\instret[31]~q ),
	.prn(vcc));
defparam \instret[31] .is_wysiwyg = "true";
defparam \instret[31] .power_up = "low";

cyclone10lp_lcell_comb \_T_198~0 (
	.dataa(\instret[0]~q ),
	.datab(\instret[1]~q ),
	.datac(\instret[31]~q ),
	.datad(\instret[30]~q ),
	.cin(gnd),
	.combout(\_T_198~0_combout ),
	.cout());
defparam \_T_198~0 .lut_mask = 16'h7FFF;
defparam \_T_198~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_198~1 (
	.dataa(\instret[29]~q ),
	.datab(\instret[28]~q ),
	.datac(\instret[27]~q ),
	.datad(\instret[26]~q ),
	.cin(gnd),
	.combout(\_T_198~1_combout ),
	.cout());
defparam \_T_198~1 .lut_mask = 16'h7FFF;
defparam \_T_198~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_198~2 (
	.dataa(\instret[25]~q ),
	.datab(\instret[24]~q ),
	.datac(\instret[23]~q ),
	.datad(\instret[22]~q ),
	.cin(gnd),
	.combout(\_T_198~2_combout ),
	.cout());
defparam \_T_198~2 .lut_mask = 16'h7FFF;
defparam \_T_198~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_198~3 (
	.dataa(\instret[21]~q ),
	.datab(\instret[20]~q ),
	.datac(\instret[19]~q ),
	.datad(\instret[18]~q ),
	.cin(gnd),
	.combout(\_T_198~3_combout ),
	.cout());
defparam \_T_198~3 .lut_mask = 16'h7FFF;
defparam \_T_198~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_198~4 (
	.dataa(\_T_198~0_combout ),
	.datab(\_T_198~1_combout ),
	.datac(\_T_198~2_combout ),
	.datad(\_T_198~3_combout ),
	.cin(gnd),
	.combout(\_T_198~4_combout ),
	.cout());
defparam \_T_198~4 .lut_mask = 16'hFFFE;
defparam \_T_198~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_198~5 (
	.dataa(\instret[17]~q ),
	.datab(\instret[16]~q ),
	.datac(\instret[15]~q ),
	.datad(\instret[14]~q ),
	.cin(gnd),
	.combout(\_T_198~5_combout ),
	.cout());
defparam \_T_198~5 .lut_mask = 16'h7FFF;
defparam \_T_198~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_198~6 (
	.dataa(\instret[13]~q ),
	.datab(\instret[12]~q ),
	.datac(\instret[11]~q ),
	.datad(\instret[10]~q ),
	.cin(gnd),
	.combout(\_T_198~6_combout ),
	.cout());
defparam \_T_198~6 .lut_mask = 16'h7FFF;
defparam \_T_198~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_198~7 (
	.dataa(\instret[9]~q ),
	.datab(\instret[8]~q ),
	.datac(\instret[7]~q ),
	.datad(\instret[6]~q ),
	.cin(gnd),
	.combout(\_T_198~7_combout ),
	.cout());
defparam \_T_198~7 .lut_mask = 16'h7FFF;
defparam \_T_198~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_198~8 (
	.dataa(\instret[5]~q ),
	.datab(\instret[4]~q ),
	.datac(\instret[3]~q ),
	.datad(\instret[2]~q ),
	.cin(gnd),
	.combout(\_T_198~8_combout ),
	.cout());
defparam \_T_198~8 .lut_mask = 16'h7FFF;
defparam \_T_198~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \_T_198~9 (
	.dataa(\_T_198~5_combout ),
	.datab(\_T_198~6_combout ),
	.datac(\_T_198~7_combout ),
	.datad(\_T_198~8_combout ),
	.cin(gnd),
	.combout(\_T_198~9_combout ),
	.cout());
defparam \_T_198~9 .lut_mask = 16'hFFFE;
defparam \_T_198~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb _T_198(
	.dataa(\isInstRet~combout ),
	.datab(\_T_198~4_combout ),
	.datac(\_T_198~9_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\_T_198~combout ),
	.cout());
defparam _T_198.lut_mask = 16'hFEFE;
defparam _T_198.sum_lutc_input = "datac";

cyclone10lp_lcell_comb \instreth[3]~38 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_198~combout ),
	.datac(gnd),
	.datad(\instreth~37_combout ),
	.cin(gnd),
	.combout(\instreth[3]~38_combout ),
	.cout());
defparam \instreth[3]~38 .lut_mask = 16'hFF77;
defparam \instreth[3]~38 .sum_lutc_input = "datac";

dffeas \instreth[0] (
	.clk(clock),
	.d(\instreth[0]~33_combout ),
	.asdata(\_T_246[0]~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[0]~q ),
	.prn(vcc));
defparam \instreth[0] .is_wysiwyg = "true";
defparam \instreth[0] .power_up = "low";

cyclone10lp_lcell_comb \instreth[1]~35 (
	.dataa(\instreth[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[0]~34 ),
	.combout(\instreth[1]~35_combout ),
	.cout(\instreth[1]~36 ));
defparam \instreth[1]~35 .lut_mask = 16'h5A5F;
defparam \instreth[1]~35 .sum_lutc_input = "cin";

dffeas \instreth[1] (
	.clk(clock),
	.d(\instreth[1]~35_combout ),
	.asdata(\_T_246[1]~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[1]~q ),
	.prn(vcc));
defparam \instreth[1] .is_wysiwyg = "true";
defparam \instreth[1] .power_up = "low";

cyclone10lp_lcell_comb \io_out[1]~15 (
	.dataa(\io_out[1]~13_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[1]~15_combout ),
	.cout());
defparam \io_out[1]~15 .lut_mask = 16'hEAEA;
defparam \io_out[1]~15 .sum_lutc_input = "datac";

dffeas \mscratch[0] (
	.clk(clock),
	.d(\_T_246[0]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[0]~q ),
	.prn(vcc));
defparam \mscratch[0] .is_wysiwyg = "true";
defparam \mscratch[0] .power_up = "low";

cyclone10lp_lcell_comb \io_out[0]~17 (
	.dataa(\mscratch[0]~q ),
	.datab(\io_out[1]~4_combout ),
	.datac(\time_[0]~q ),
	.datad(\Equal25~3_combout ),
	.cin(gnd),
	.combout(\io_out[0]~17_combout ),
	.cout());
defparam \io_out[0]~17 .lut_mask = 16'hEAC0;
defparam \io_out[0]~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[0]~18 (
	.dataa(mepc_0),
	.datab(\io_out[1]~12_combout ),
	.datac(\timeh[0]~q ),
	.datad(\Equal26~0_combout ),
	.cin(gnd),
	.combout(\io_out[0]~18_combout ),
	.cout());
defparam \io_out[0]~18 .lut_mask = 16'hEAC0;
defparam \io_out[0]~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mcause[0]~12 (
	.dataa(isEcall),
	.datab(io_expt1),
	.datac(\_T_246[0]~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mcause[0]~12_combout ),
	.cout());
defparam \mcause[0]~12 .lut_mask = 16'hEAEA;
defparam \mcause[0]~12 .sum_lutc_input = "datac";

dffeas \mcause[0] (
	.clk(clock),
	.d(\mcause[0]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mcause[0]~11_combout ),
	.q(\mcause[0]~q ),
	.prn(vcc));
defparam \mcause[0] .is_wysiwyg = "true";
defparam \mcause[0] .power_up = "low";

cyclone10lp_lcell_comb \io_out[0]~19 (
	.dataa(\mcause[0]~q ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[0]~q ),
	.datad(\Equal27~0_combout ),
	.cin(gnd),
	.combout(\io_out[0]~19_combout ),
	.cout());
defparam \io_out[0]~19 .lut_mask = 16'hEAC0;
defparam \io_out[0]~19 .sum_lutc_input = "datac";

dffeas \mbadaddr[0] (
	.clk(clock),
	.d(\_T_246[0]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[0]~q ),
	.prn(vcc));
defparam \mbadaddr[0] .is_wysiwyg = "true";
defparam \mbadaddr[0] .power_up = "low";

cyclone10lp_lcell_comb \io_out[0]~20 (
	.dataa(\mbadaddr[0]~q ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[0]~q ),
	.datad(\Equal28~0_combout ),
	.cin(gnd),
	.combout(\io_out[0]~20_combout ),
	.cout());
defparam \io_out[0]~20 .lut_mask = 16'hEAC0;
defparam \io_out[0]~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[0]~21 (
	.dataa(\io_out[0]~17_combout ),
	.datab(\io_out[0]~18_combout ),
	.datac(\io_out[0]~19_combout ),
	.datad(\io_out[0]~20_combout ),
	.cin(gnd),
	.combout(\io_out[0]~21_combout ),
	.cout());
defparam \io_out[0]~21 .lut_mask = 16'hFFFE;
defparam \io_out[0]~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \IE~2 (
	.dataa(io_expt1),
	.datab(isEcall),
	.datac(altera_reset_synchronizer_int_chain_out),
	.datad(\_T_246[0]~2_combout ),
	.cin(gnd),
	.combout(\IE~2_combout ),
	.cout());
defparam \IE~2 .lut_mask = 16'h2000;
defparam \IE~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \IE1~0 (
	.dataa(io_expt2),
	.datab(\Equal30~0_combout ),
	.datac(\wen~combout ),
	.datad(mcause_0),
	.cin(gnd),
	.combout(\IE1~0_combout ),
	.cout());
defparam \IE1~0 .lut_mask = 16'h2AFF;
defparam \IE1~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \PRV1[0]~4 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\IE1~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\PRV1[0]~4_combout ),
	.cout());
defparam \PRV1[0]~4 .lut_mask = 16'h7777;
defparam \PRV1[0]~4 .sum_lutc_input = "datac";

dffeas IE(
	.clk(clock),
	.d(\IE~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PRV1[0]~4_combout ),
	.q(\IE~q ),
	.prn(vcc));
defparam IE.is_wysiwyg = "true";
defparam IE.power_up = "low";

cyclone10lp_lcell_comb \io_out[0]~22 (
	.dataa(mtvec_0),
	.datab(\IE~q ),
	.datac(\Equal30~0_combout ),
	.datad(\Equal19~3_combout ),
	.cin(gnd),
	.combout(\io_out[0]~22_combout ),
	.cout());
defparam \io_out[0]~22 .lut_mask = 16'hEAC0;
defparam \io_out[0]~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[0]~23 (
	.dataa(\io_out[0]~22_combout ),
	.datab(\io_out[1]~10_combout ),
	.datac(\cycleh[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[0]~23_combout ),
	.cout());
defparam \io_out[0]~23 .lut_mask = 16'hEAEA;
defparam \io_out[0]~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_246[2]~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~3_combout ),
	.cout());
defparam \mtvec~3 .lut_mask = 16'h8888;
defparam \mtvec~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~4 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_246[3]~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~4_combout ),
	.cout());
defparam \mtvec~4 .lut_mask = 16'h8888;
defparam \mtvec~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~5 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[4]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~5_combout ),
	.cout());
defparam \mtvec~5 .lut_mask = 16'h8888;
defparam \mtvec~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~6 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[5]~3_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~6_combout ),
	.cout());
defparam \mtvec~6 .lut_mask = 16'h8888;
defparam \mtvec~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~7 (
	.dataa(\_T_244[6]~5_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\mtvec~7_combout ),
	.cout());
defparam \mtvec~7 .lut_mask = 16'hAAFF;
defparam \mtvec~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~8 (
	.dataa(\_T_244[7]~7_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\mtvec~8_combout ),
	.cout());
defparam \mtvec~8 .lut_mask = 16'hAAFF;
defparam \mtvec~8 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~9 (
	.dataa(\_T_244[8]~9_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\mtvec~9_combout ),
	.cout());
defparam \mtvec~9 .lut_mask = 16'hAAFF;
defparam \mtvec~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~10 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[9]~11_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~10_combout ),
	.cout());
defparam \mtvec~10 .lut_mask = 16'h8888;
defparam \mtvec~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~11 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[10]~13_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~11_combout ),
	.cout());
defparam \mtvec~11 .lut_mask = 16'h8888;
defparam \mtvec~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~12 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[11]~15_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~12_combout ),
	.cout());
defparam \mtvec~12 .lut_mask = 16'h8888;
defparam \mtvec~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~13 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[12]~17_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~13_combout ),
	.cout());
defparam \mtvec~13 .lut_mask = 16'h8888;
defparam \mtvec~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~14 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[13]~19_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~14_combout ),
	.cout());
defparam \mtvec~14 .lut_mask = 16'h8888;
defparam \mtvec~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~15 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[14]~21_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~15_combout ),
	.cout());
defparam \mtvec~15 .lut_mask = 16'h8888;
defparam \mtvec~15 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~16 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[15]~23_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~16_combout ),
	.cout());
defparam \mtvec~16 .lut_mask = 16'h8888;
defparam \mtvec~16 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~17 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[16]~25_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~17_combout ),
	.cout());
defparam \mtvec~17 .lut_mask = 16'h8888;
defparam \mtvec~17 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~18 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[17]~27_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~18_combout ),
	.cout());
defparam \mtvec~18 .lut_mask = 16'h8888;
defparam \mtvec~18 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~19 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[18]~29_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~19_combout ),
	.cout());
defparam \mtvec~19 .lut_mask = 16'h8888;
defparam \mtvec~19 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~20 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[19]~31_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~20_combout ),
	.cout());
defparam \mtvec~20 .lut_mask = 16'h8888;
defparam \mtvec~20 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~21 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[20]~33_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~21_combout ),
	.cout());
defparam \mtvec~21 .lut_mask = 16'h8888;
defparam \mtvec~21 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~22 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[21]~35_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~22_combout ),
	.cout());
defparam \mtvec~22 .lut_mask = 16'h8888;
defparam \mtvec~22 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~23 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[22]~37_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~23_combout ),
	.cout());
defparam \mtvec~23 .lut_mask = 16'h8888;
defparam \mtvec~23 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~24 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[23]~39_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~24_combout ),
	.cout());
defparam \mtvec~24 .lut_mask = 16'h8888;
defparam \mtvec~24 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~25 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[24]~41_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~25_combout ),
	.cout());
defparam \mtvec~25 .lut_mask = 16'h8888;
defparam \mtvec~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~26 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[25]~43_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~26_combout ),
	.cout());
defparam \mtvec~26 .lut_mask = 16'h8888;
defparam \mtvec~26 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~27 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[26]~45_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~27_combout ),
	.cout());
defparam \mtvec~27 .lut_mask = 16'h8888;
defparam \mtvec~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~28 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[27]~47_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~28_combout ),
	.cout());
defparam \mtvec~28 .lut_mask = 16'h8888;
defparam \mtvec~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~29 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[28]~49_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~29_combout ),
	.cout());
defparam \mtvec~29 .lut_mask = 16'h8888;
defparam \mtvec~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~30 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[29]~51_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~30_combout ),
	.cout());
defparam \mtvec~30 .lut_mask = 16'h8888;
defparam \mtvec~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~31 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[30]~53_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~31_combout ),
	.cout());
defparam \mtvec~31 .lut_mask = 16'h8888;
defparam \mtvec~31 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mtvec~32 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_246[31]~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mtvec~32_combout ),
	.cout());
defparam \mtvec~32 .lut_mask = 16'h8888;
defparam \mtvec~32 .sum_lutc_input = "datac";

dffeas \mscratch[28] (
	.clk(clock),
	.d(\_T_244[28]~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[28]~q ),
	.prn(vcc));
defparam \mscratch[28] .is_wysiwyg = "true";
defparam \mscratch[28] .power_up = "low";

cyclone10lp_lcell_comb \io_out[28]~25 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[28]~q ),
	.datad(\mscratch[28]~q ),
	.cin(gnd),
	.combout(\io_out[28]~25_combout ),
	.cout());
defparam \io_out[28]~25 .lut_mask = 16'hEAC0;
defparam \io_out[28]~25 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[28]~26 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_28),
	.datad(\time_[28]~q ),
	.cin(gnd),
	.combout(\io_out[28]~26_combout ),
	.cout());
defparam \io_out[28]~26 .lut_mask = 16'hEAC0;
defparam \io_out[28]~26 .sum_lutc_input = "datac";

dffeas \mbadaddr[28] (
	.clk(clock),
	.d(\_T_244[28]~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[28]~q ),
	.prn(vcc));
defparam \mbadaddr[28] .is_wysiwyg = "true";
defparam \mbadaddr[28] .power_up = "low";

cyclone10lp_lcell_comb \io_out[28]~27 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[28]~q ),
	.datad(\mbadaddr[28]~q ),
	.cin(gnd),
	.combout(\io_out[28]~27_combout ),
	.cout());
defparam \io_out[28]~27 .lut_mask = 16'hEAC0;
defparam \io_out[28]~27 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cycleh[2]~38 (
	.dataa(\cycleh[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[1]~35 ),
	.combout(\cycleh[2]~38_combout ),
	.cout(\cycleh[2]~39 ));
defparam \cycleh[2]~38 .lut_mask = 16'hA50A;
defparam \cycleh[2]~38 .sum_lutc_input = "cin";

dffeas \cycleh[2] (
	.clk(clock),
	.d(\cycleh[2]~38_combout ),
	.asdata(\_T_246[2]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[2]~q ),
	.prn(vcc));
defparam \cycleh[2] .is_wysiwyg = "true";
defparam \cycleh[2] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[3]~40 (
	.dataa(\cycleh[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[2]~39 ),
	.combout(\cycleh[3]~40_combout ),
	.cout(\cycleh[3]~41 ));
defparam \cycleh[3]~40 .lut_mask = 16'h5A5F;
defparam \cycleh[3]~40 .sum_lutc_input = "cin";

dffeas \cycleh[3] (
	.clk(clock),
	.d(\cycleh[3]~40_combout ),
	.asdata(\_T_246[3]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[3]~q ),
	.prn(vcc));
defparam \cycleh[3] .is_wysiwyg = "true";
defparam \cycleh[3] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[4]~42 (
	.dataa(\cycleh[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[3]~41 ),
	.combout(\cycleh[4]~42_combout ),
	.cout(\cycleh[4]~43 ));
defparam \cycleh[4]~42 .lut_mask = 16'hA50A;
defparam \cycleh[4]~42 .sum_lutc_input = "cin";

dffeas \cycleh[4] (
	.clk(clock),
	.d(\cycleh[4]~42_combout ),
	.asdata(\_T_244[4]~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[4]~q ),
	.prn(vcc));
defparam \cycleh[4] .is_wysiwyg = "true";
defparam \cycleh[4] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[5]~44 (
	.dataa(\cycleh[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[4]~43 ),
	.combout(\cycleh[5]~44_combout ),
	.cout(\cycleh[5]~45 ));
defparam \cycleh[5]~44 .lut_mask = 16'h5A5F;
defparam \cycleh[5]~44 .sum_lutc_input = "cin";

dffeas \cycleh[5] (
	.clk(clock),
	.d(\cycleh[5]~44_combout ),
	.asdata(\_T_244[5]~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[5]~q ),
	.prn(vcc));
defparam \cycleh[5] .is_wysiwyg = "true";
defparam \cycleh[5] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[6]~46 (
	.dataa(\cycleh[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[5]~45 ),
	.combout(\cycleh[6]~46_combout ),
	.cout(\cycleh[6]~47 ));
defparam \cycleh[6]~46 .lut_mask = 16'hA50A;
defparam \cycleh[6]~46 .sum_lutc_input = "cin";

dffeas \cycleh[6] (
	.clk(clock),
	.d(\cycleh[6]~46_combout ),
	.asdata(\_T_244[6]~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[6]~q ),
	.prn(vcc));
defparam \cycleh[6] .is_wysiwyg = "true";
defparam \cycleh[6] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[7]~48 (
	.dataa(\cycleh[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[6]~47 ),
	.combout(\cycleh[7]~48_combout ),
	.cout(\cycleh[7]~49 ));
defparam \cycleh[7]~48 .lut_mask = 16'h5A5F;
defparam \cycleh[7]~48 .sum_lutc_input = "cin";

dffeas \cycleh[7] (
	.clk(clock),
	.d(\cycleh[7]~48_combout ),
	.asdata(\_T_244[7]~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[7]~q ),
	.prn(vcc));
defparam \cycleh[7] .is_wysiwyg = "true";
defparam \cycleh[7] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[8]~50 (
	.dataa(\cycleh[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[7]~49 ),
	.combout(\cycleh[8]~50_combout ),
	.cout(\cycleh[8]~51 ));
defparam \cycleh[8]~50 .lut_mask = 16'hA50A;
defparam \cycleh[8]~50 .sum_lutc_input = "cin";

dffeas \cycleh[8] (
	.clk(clock),
	.d(\cycleh[8]~50_combout ),
	.asdata(\_T_244[8]~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[8]~q ),
	.prn(vcc));
defparam \cycleh[8] .is_wysiwyg = "true";
defparam \cycleh[8] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[9]~52 (
	.dataa(\cycleh[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[8]~51 ),
	.combout(\cycleh[9]~52_combout ),
	.cout(\cycleh[9]~53 ));
defparam \cycleh[9]~52 .lut_mask = 16'h5A5F;
defparam \cycleh[9]~52 .sum_lutc_input = "cin";

dffeas \cycleh[9] (
	.clk(clock),
	.d(\cycleh[9]~52_combout ),
	.asdata(\_T_244[9]~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[9]~q ),
	.prn(vcc));
defparam \cycleh[9] .is_wysiwyg = "true";
defparam \cycleh[9] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[10]~54 (
	.dataa(\cycleh[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[9]~53 ),
	.combout(\cycleh[10]~54_combout ),
	.cout(\cycleh[10]~55 ));
defparam \cycleh[10]~54 .lut_mask = 16'hA50A;
defparam \cycleh[10]~54 .sum_lutc_input = "cin";

dffeas \cycleh[10] (
	.clk(clock),
	.d(\cycleh[10]~54_combout ),
	.asdata(\_T_244[10]~13_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[10]~q ),
	.prn(vcc));
defparam \cycleh[10] .is_wysiwyg = "true";
defparam \cycleh[10] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[11]~56 (
	.dataa(\cycleh[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[10]~55 ),
	.combout(\cycleh[11]~56_combout ),
	.cout(\cycleh[11]~57 ));
defparam \cycleh[11]~56 .lut_mask = 16'h5A5F;
defparam \cycleh[11]~56 .sum_lutc_input = "cin";

dffeas \cycleh[11] (
	.clk(clock),
	.d(\cycleh[11]~56_combout ),
	.asdata(\_T_244[11]~15_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[11]~q ),
	.prn(vcc));
defparam \cycleh[11] .is_wysiwyg = "true";
defparam \cycleh[11] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[12]~58 (
	.dataa(\cycleh[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[11]~57 ),
	.combout(\cycleh[12]~58_combout ),
	.cout(\cycleh[12]~59 ));
defparam \cycleh[12]~58 .lut_mask = 16'hA50A;
defparam \cycleh[12]~58 .sum_lutc_input = "cin";

dffeas \cycleh[12] (
	.clk(clock),
	.d(\cycleh[12]~58_combout ),
	.asdata(\_T_244[12]~17_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[12]~q ),
	.prn(vcc));
defparam \cycleh[12] .is_wysiwyg = "true";
defparam \cycleh[12] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[13]~60 (
	.dataa(\cycleh[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[12]~59 ),
	.combout(\cycleh[13]~60_combout ),
	.cout(\cycleh[13]~61 ));
defparam \cycleh[13]~60 .lut_mask = 16'h5A5F;
defparam \cycleh[13]~60 .sum_lutc_input = "cin";

dffeas \cycleh[13] (
	.clk(clock),
	.d(\cycleh[13]~60_combout ),
	.asdata(\_T_244[13]~19_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[13]~q ),
	.prn(vcc));
defparam \cycleh[13] .is_wysiwyg = "true";
defparam \cycleh[13] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[14]~62 (
	.dataa(\cycleh[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[13]~61 ),
	.combout(\cycleh[14]~62_combout ),
	.cout(\cycleh[14]~63 ));
defparam \cycleh[14]~62 .lut_mask = 16'hA50A;
defparam \cycleh[14]~62 .sum_lutc_input = "cin";

dffeas \cycleh[14] (
	.clk(clock),
	.d(\cycleh[14]~62_combout ),
	.asdata(\_T_244[14]~21_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[14]~q ),
	.prn(vcc));
defparam \cycleh[14] .is_wysiwyg = "true";
defparam \cycleh[14] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[15]~64 (
	.dataa(\cycleh[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[14]~63 ),
	.combout(\cycleh[15]~64_combout ),
	.cout(\cycleh[15]~65 ));
defparam \cycleh[15]~64 .lut_mask = 16'h5A5F;
defparam \cycleh[15]~64 .sum_lutc_input = "cin";

dffeas \cycleh[15] (
	.clk(clock),
	.d(\cycleh[15]~64_combout ),
	.asdata(\_T_244[15]~23_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[15]~q ),
	.prn(vcc));
defparam \cycleh[15] .is_wysiwyg = "true";
defparam \cycleh[15] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[16]~66 (
	.dataa(\cycleh[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[15]~65 ),
	.combout(\cycleh[16]~66_combout ),
	.cout(\cycleh[16]~67 ));
defparam \cycleh[16]~66 .lut_mask = 16'hA50A;
defparam \cycleh[16]~66 .sum_lutc_input = "cin";

dffeas \cycleh[16] (
	.clk(clock),
	.d(\cycleh[16]~66_combout ),
	.asdata(\_T_244[16]~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[16]~q ),
	.prn(vcc));
defparam \cycleh[16] .is_wysiwyg = "true";
defparam \cycleh[16] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[17]~68 (
	.dataa(\cycleh[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[16]~67 ),
	.combout(\cycleh[17]~68_combout ),
	.cout(\cycleh[17]~69 ));
defparam \cycleh[17]~68 .lut_mask = 16'h5A5F;
defparam \cycleh[17]~68 .sum_lutc_input = "cin";

dffeas \cycleh[17] (
	.clk(clock),
	.d(\cycleh[17]~68_combout ),
	.asdata(\_T_244[17]~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[17]~q ),
	.prn(vcc));
defparam \cycleh[17] .is_wysiwyg = "true";
defparam \cycleh[17] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[18]~70 (
	.dataa(\cycleh[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[17]~69 ),
	.combout(\cycleh[18]~70_combout ),
	.cout(\cycleh[18]~71 ));
defparam \cycleh[18]~70 .lut_mask = 16'hA50A;
defparam \cycleh[18]~70 .sum_lutc_input = "cin";

dffeas \cycleh[18] (
	.clk(clock),
	.d(\cycleh[18]~70_combout ),
	.asdata(\_T_244[18]~29_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[18]~q ),
	.prn(vcc));
defparam \cycleh[18] .is_wysiwyg = "true";
defparam \cycleh[18] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[19]~72 (
	.dataa(\cycleh[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[18]~71 ),
	.combout(\cycleh[19]~72_combout ),
	.cout(\cycleh[19]~73 ));
defparam \cycleh[19]~72 .lut_mask = 16'h5A5F;
defparam \cycleh[19]~72 .sum_lutc_input = "cin";

dffeas \cycleh[19] (
	.clk(clock),
	.d(\cycleh[19]~72_combout ),
	.asdata(\_T_244[19]~31_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[19]~q ),
	.prn(vcc));
defparam \cycleh[19] .is_wysiwyg = "true";
defparam \cycleh[19] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[20]~74 (
	.dataa(\cycleh[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[19]~73 ),
	.combout(\cycleh[20]~74_combout ),
	.cout(\cycleh[20]~75 ));
defparam \cycleh[20]~74 .lut_mask = 16'hA50A;
defparam \cycleh[20]~74 .sum_lutc_input = "cin";

dffeas \cycleh[20] (
	.clk(clock),
	.d(\cycleh[20]~74_combout ),
	.asdata(\_T_244[20]~33_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[20]~q ),
	.prn(vcc));
defparam \cycleh[20] .is_wysiwyg = "true";
defparam \cycleh[20] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[21]~76 (
	.dataa(\cycleh[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[20]~75 ),
	.combout(\cycleh[21]~76_combout ),
	.cout(\cycleh[21]~77 ));
defparam \cycleh[21]~76 .lut_mask = 16'h5A5F;
defparam \cycleh[21]~76 .sum_lutc_input = "cin";

dffeas \cycleh[21] (
	.clk(clock),
	.d(\cycleh[21]~76_combout ),
	.asdata(\_T_244[21]~35_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[21]~q ),
	.prn(vcc));
defparam \cycleh[21] .is_wysiwyg = "true";
defparam \cycleh[21] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[22]~78 (
	.dataa(\cycleh[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[21]~77 ),
	.combout(\cycleh[22]~78_combout ),
	.cout(\cycleh[22]~79 ));
defparam \cycleh[22]~78 .lut_mask = 16'hA50A;
defparam \cycleh[22]~78 .sum_lutc_input = "cin";

dffeas \cycleh[22] (
	.clk(clock),
	.d(\cycleh[22]~78_combout ),
	.asdata(\_T_244[22]~37_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[22]~q ),
	.prn(vcc));
defparam \cycleh[22] .is_wysiwyg = "true";
defparam \cycleh[22] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[23]~80 (
	.dataa(\cycleh[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[22]~79 ),
	.combout(\cycleh[23]~80_combout ),
	.cout(\cycleh[23]~81 ));
defparam \cycleh[23]~80 .lut_mask = 16'h5A5F;
defparam \cycleh[23]~80 .sum_lutc_input = "cin";

dffeas \cycleh[23] (
	.clk(clock),
	.d(\cycleh[23]~80_combout ),
	.asdata(\_T_244[23]~39_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[23]~q ),
	.prn(vcc));
defparam \cycleh[23] .is_wysiwyg = "true";
defparam \cycleh[23] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[24]~82 (
	.dataa(\cycleh[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[23]~81 ),
	.combout(\cycleh[24]~82_combout ),
	.cout(\cycleh[24]~83 ));
defparam \cycleh[24]~82 .lut_mask = 16'hA50A;
defparam \cycleh[24]~82 .sum_lutc_input = "cin";

dffeas \cycleh[24] (
	.clk(clock),
	.d(\cycleh[24]~82_combout ),
	.asdata(\_T_244[24]~41_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[24]~q ),
	.prn(vcc));
defparam \cycleh[24] .is_wysiwyg = "true";
defparam \cycleh[24] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[25]~84 (
	.dataa(\cycleh[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[24]~83 ),
	.combout(\cycleh[25]~84_combout ),
	.cout(\cycleh[25]~85 ));
defparam \cycleh[25]~84 .lut_mask = 16'h5A5F;
defparam \cycleh[25]~84 .sum_lutc_input = "cin";

dffeas \cycleh[25] (
	.clk(clock),
	.d(\cycleh[25]~84_combout ),
	.asdata(\_T_244[25]~43_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[25]~q ),
	.prn(vcc));
defparam \cycleh[25] .is_wysiwyg = "true";
defparam \cycleh[25] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[26]~86 (
	.dataa(\cycleh[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[25]~85 ),
	.combout(\cycleh[26]~86_combout ),
	.cout(\cycleh[26]~87 ));
defparam \cycleh[26]~86 .lut_mask = 16'hA50A;
defparam \cycleh[26]~86 .sum_lutc_input = "cin";

dffeas \cycleh[26] (
	.clk(clock),
	.d(\cycleh[26]~86_combout ),
	.asdata(\_T_244[26]~45_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[26]~q ),
	.prn(vcc));
defparam \cycleh[26] .is_wysiwyg = "true";
defparam \cycleh[26] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[27]~88 (
	.dataa(\cycleh[27]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[26]~87 ),
	.combout(\cycleh[27]~88_combout ),
	.cout(\cycleh[27]~89 ));
defparam \cycleh[27]~88 .lut_mask = 16'h5A5F;
defparam \cycleh[27]~88 .sum_lutc_input = "cin";

dffeas \cycleh[27] (
	.clk(clock),
	.d(\cycleh[27]~88_combout ),
	.asdata(\_T_244[27]~47_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[27]~q ),
	.prn(vcc));
defparam \cycleh[27] .is_wysiwyg = "true";
defparam \cycleh[27] .power_up = "low";

cyclone10lp_lcell_comb \cycleh[28]~90 (
	.dataa(\cycleh[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[27]~89 ),
	.combout(\cycleh[28]~90_combout ),
	.cout(\cycleh[28]~91 ));
defparam \cycleh[28]~90 .lut_mask = 16'hA50A;
defparam \cycleh[28]~90 .sum_lutc_input = "cin";

dffeas \cycleh[28] (
	.clk(clock),
	.d(\cycleh[28]~90_combout ),
	.asdata(\_T_244[28]~49_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[28]~q ),
	.prn(vcc));
defparam \cycleh[28] .is_wysiwyg = "true";
defparam \cycleh[28] .power_up = "low";

cyclone10lp_lcell_comb \io_out[28]~28 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_28),
	.datad(\cycleh[28]~q ),
	.cin(gnd),
	.combout(\io_out[28]~28_combout ),
	.cout());
defparam \io_out[28]~28 .lut_mask = 16'hEAC0;
defparam \io_out[28]~28 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[28]~29 (
	.dataa(\io_out[28]~25_combout ),
	.datab(\io_out[28]~26_combout ),
	.datac(\io_out[28]~27_combout ),
	.datad(\io_out[28]~28_combout ),
	.cin(gnd),
	.combout(\io_out[28]~29_combout ),
	.cout());
defparam \io_out[28]~29 .lut_mask = 16'hFFFE;
defparam \io_out[28]~29 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \instreth[2]~39 (
	.dataa(\instreth[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[1]~36 ),
	.combout(\instreth[2]~39_combout ),
	.cout(\instreth[2]~40 ));
defparam \instreth[2]~39 .lut_mask = 16'hA50A;
defparam \instreth[2]~39 .sum_lutc_input = "cin";

dffeas \instreth[2] (
	.clk(clock),
	.d(\instreth[2]~39_combout ),
	.asdata(\_T_246[2]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[2]~q ),
	.prn(vcc));
defparam \instreth[2] .is_wysiwyg = "true";
defparam \instreth[2] .power_up = "low";

cyclone10lp_lcell_comb \instreth[3]~41 (
	.dataa(\instreth[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[2]~40 ),
	.combout(\instreth[3]~41_combout ),
	.cout(\instreth[3]~42 ));
defparam \instreth[3]~41 .lut_mask = 16'h5A5F;
defparam \instreth[3]~41 .sum_lutc_input = "cin";

dffeas \instreth[3] (
	.clk(clock),
	.d(\instreth[3]~41_combout ),
	.asdata(\_T_246[3]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[3]~q ),
	.prn(vcc));
defparam \instreth[3] .is_wysiwyg = "true";
defparam \instreth[3] .power_up = "low";

cyclone10lp_lcell_comb \instreth[4]~43 (
	.dataa(\instreth[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[3]~42 ),
	.combout(\instreth[4]~43_combout ),
	.cout(\instreth[4]~44 ));
defparam \instreth[4]~43 .lut_mask = 16'hA50A;
defparam \instreth[4]~43 .sum_lutc_input = "cin";

dffeas \instreth[4] (
	.clk(clock),
	.d(\instreth[4]~43_combout ),
	.asdata(\_T_244[4]~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[4]~q ),
	.prn(vcc));
defparam \instreth[4] .is_wysiwyg = "true";
defparam \instreth[4] .power_up = "low";

cyclone10lp_lcell_comb \instreth[5]~45 (
	.dataa(\instreth[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[4]~44 ),
	.combout(\instreth[5]~45_combout ),
	.cout(\instreth[5]~46 ));
defparam \instreth[5]~45 .lut_mask = 16'h5A5F;
defparam \instreth[5]~45 .sum_lutc_input = "cin";

dffeas \instreth[5] (
	.clk(clock),
	.d(\instreth[5]~45_combout ),
	.asdata(\_T_244[5]~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[5]~q ),
	.prn(vcc));
defparam \instreth[5] .is_wysiwyg = "true";
defparam \instreth[5] .power_up = "low";

cyclone10lp_lcell_comb \instreth[6]~47 (
	.dataa(\instreth[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[5]~46 ),
	.combout(\instreth[6]~47_combout ),
	.cout(\instreth[6]~48 ));
defparam \instreth[6]~47 .lut_mask = 16'hA50A;
defparam \instreth[6]~47 .sum_lutc_input = "cin";

dffeas \instreth[6] (
	.clk(clock),
	.d(\instreth[6]~47_combout ),
	.asdata(\_T_244[6]~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[6]~q ),
	.prn(vcc));
defparam \instreth[6] .is_wysiwyg = "true";
defparam \instreth[6] .power_up = "low";

cyclone10lp_lcell_comb \instreth[7]~49 (
	.dataa(\instreth[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[6]~48 ),
	.combout(\instreth[7]~49_combout ),
	.cout(\instreth[7]~50 ));
defparam \instreth[7]~49 .lut_mask = 16'h5A5F;
defparam \instreth[7]~49 .sum_lutc_input = "cin";

dffeas \instreth[7] (
	.clk(clock),
	.d(\instreth[7]~49_combout ),
	.asdata(\_T_244[7]~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[7]~q ),
	.prn(vcc));
defparam \instreth[7] .is_wysiwyg = "true";
defparam \instreth[7] .power_up = "low";

cyclone10lp_lcell_comb \instreth[8]~51 (
	.dataa(\instreth[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[7]~50 ),
	.combout(\instreth[8]~51_combout ),
	.cout(\instreth[8]~52 ));
defparam \instreth[8]~51 .lut_mask = 16'hA50A;
defparam \instreth[8]~51 .sum_lutc_input = "cin";

dffeas \instreth[8] (
	.clk(clock),
	.d(\instreth[8]~51_combout ),
	.asdata(\_T_244[8]~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[8]~q ),
	.prn(vcc));
defparam \instreth[8] .is_wysiwyg = "true";
defparam \instreth[8] .power_up = "low";

cyclone10lp_lcell_comb \instreth[9]~53 (
	.dataa(\instreth[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[8]~52 ),
	.combout(\instreth[9]~53_combout ),
	.cout(\instreth[9]~54 ));
defparam \instreth[9]~53 .lut_mask = 16'h5A5F;
defparam \instreth[9]~53 .sum_lutc_input = "cin";

dffeas \instreth[9] (
	.clk(clock),
	.d(\instreth[9]~53_combout ),
	.asdata(\_T_244[9]~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[9]~q ),
	.prn(vcc));
defparam \instreth[9] .is_wysiwyg = "true";
defparam \instreth[9] .power_up = "low";

cyclone10lp_lcell_comb \instreth[10]~55 (
	.dataa(\instreth[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[9]~54 ),
	.combout(\instreth[10]~55_combout ),
	.cout(\instreth[10]~56 ));
defparam \instreth[10]~55 .lut_mask = 16'hA50A;
defparam \instreth[10]~55 .sum_lutc_input = "cin";

dffeas \instreth[10] (
	.clk(clock),
	.d(\instreth[10]~55_combout ),
	.asdata(\_T_244[10]~13_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[10]~q ),
	.prn(vcc));
defparam \instreth[10] .is_wysiwyg = "true";
defparam \instreth[10] .power_up = "low";

cyclone10lp_lcell_comb \instreth[11]~57 (
	.dataa(\instreth[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[10]~56 ),
	.combout(\instreth[11]~57_combout ),
	.cout(\instreth[11]~58 ));
defparam \instreth[11]~57 .lut_mask = 16'h5A5F;
defparam \instreth[11]~57 .sum_lutc_input = "cin";

dffeas \instreth[11] (
	.clk(clock),
	.d(\instreth[11]~57_combout ),
	.asdata(\_T_244[11]~15_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[11]~q ),
	.prn(vcc));
defparam \instreth[11] .is_wysiwyg = "true";
defparam \instreth[11] .power_up = "low";

cyclone10lp_lcell_comb \instreth[12]~59 (
	.dataa(\instreth[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[11]~58 ),
	.combout(\instreth[12]~59_combout ),
	.cout(\instreth[12]~60 ));
defparam \instreth[12]~59 .lut_mask = 16'hA50A;
defparam \instreth[12]~59 .sum_lutc_input = "cin";

dffeas \instreth[12] (
	.clk(clock),
	.d(\instreth[12]~59_combout ),
	.asdata(\_T_244[12]~17_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[12]~q ),
	.prn(vcc));
defparam \instreth[12] .is_wysiwyg = "true";
defparam \instreth[12] .power_up = "low";

cyclone10lp_lcell_comb \instreth[13]~61 (
	.dataa(\instreth[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[12]~60 ),
	.combout(\instreth[13]~61_combout ),
	.cout(\instreth[13]~62 ));
defparam \instreth[13]~61 .lut_mask = 16'h5A5F;
defparam \instreth[13]~61 .sum_lutc_input = "cin";

dffeas \instreth[13] (
	.clk(clock),
	.d(\instreth[13]~61_combout ),
	.asdata(\_T_244[13]~19_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[13]~q ),
	.prn(vcc));
defparam \instreth[13] .is_wysiwyg = "true";
defparam \instreth[13] .power_up = "low";

cyclone10lp_lcell_comb \instreth[14]~63 (
	.dataa(\instreth[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[13]~62 ),
	.combout(\instreth[14]~63_combout ),
	.cout(\instreth[14]~64 ));
defparam \instreth[14]~63 .lut_mask = 16'hA50A;
defparam \instreth[14]~63 .sum_lutc_input = "cin";

dffeas \instreth[14] (
	.clk(clock),
	.d(\instreth[14]~63_combout ),
	.asdata(\_T_244[14]~21_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[14]~q ),
	.prn(vcc));
defparam \instreth[14] .is_wysiwyg = "true";
defparam \instreth[14] .power_up = "low";

cyclone10lp_lcell_comb \instreth[15]~65 (
	.dataa(\instreth[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[14]~64 ),
	.combout(\instreth[15]~65_combout ),
	.cout(\instreth[15]~66 ));
defparam \instreth[15]~65 .lut_mask = 16'h5A5F;
defparam \instreth[15]~65 .sum_lutc_input = "cin";

dffeas \instreth[15] (
	.clk(clock),
	.d(\instreth[15]~65_combout ),
	.asdata(\_T_244[15]~23_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[15]~q ),
	.prn(vcc));
defparam \instreth[15] .is_wysiwyg = "true";
defparam \instreth[15] .power_up = "low";

cyclone10lp_lcell_comb \instreth[16]~67 (
	.dataa(\instreth[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[15]~66 ),
	.combout(\instreth[16]~67_combout ),
	.cout(\instreth[16]~68 ));
defparam \instreth[16]~67 .lut_mask = 16'hA50A;
defparam \instreth[16]~67 .sum_lutc_input = "cin";

dffeas \instreth[16] (
	.clk(clock),
	.d(\instreth[16]~67_combout ),
	.asdata(\_T_244[16]~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[16]~q ),
	.prn(vcc));
defparam \instreth[16] .is_wysiwyg = "true";
defparam \instreth[16] .power_up = "low";

cyclone10lp_lcell_comb \instreth[17]~69 (
	.dataa(\instreth[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[16]~68 ),
	.combout(\instreth[17]~69_combout ),
	.cout(\instreth[17]~70 ));
defparam \instreth[17]~69 .lut_mask = 16'h5A5F;
defparam \instreth[17]~69 .sum_lutc_input = "cin";

dffeas \instreth[17] (
	.clk(clock),
	.d(\instreth[17]~69_combout ),
	.asdata(\_T_244[17]~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[17]~q ),
	.prn(vcc));
defparam \instreth[17] .is_wysiwyg = "true";
defparam \instreth[17] .power_up = "low";

cyclone10lp_lcell_comb \instreth[18]~71 (
	.dataa(\instreth[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[17]~70 ),
	.combout(\instreth[18]~71_combout ),
	.cout(\instreth[18]~72 ));
defparam \instreth[18]~71 .lut_mask = 16'hA50A;
defparam \instreth[18]~71 .sum_lutc_input = "cin";

dffeas \instreth[18] (
	.clk(clock),
	.d(\instreth[18]~71_combout ),
	.asdata(\_T_244[18]~29_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[18]~q ),
	.prn(vcc));
defparam \instreth[18] .is_wysiwyg = "true";
defparam \instreth[18] .power_up = "low";

cyclone10lp_lcell_comb \instreth[19]~73 (
	.dataa(\instreth[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[18]~72 ),
	.combout(\instreth[19]~73_combout ),
	.cout(\instreth[19]~74 ));
defparam \instreth[19]~73 .lut_mask = 16'h5A5F;
defparam \instreth[19]~73 .sum_lutc_input = "cin";

dffeas \instreth[19] (
	.clk(clock),
	.d(\instreth[19]~73_combout ),
	.asdata(\_T_244[19]~31_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[19]~q ),
	.prn(vcc));
defparam \instreth[19] .is_wysiwyg = "true";
defparam \instreth[19] .power_up = "low";

cyclone10lp_lcell_comb \instreth[20]~75 (
	.dataa(\instreth[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[19]~74 ),
	.combout(\instreth[20]~75_combout ),
	.cout(\instreth[20]~76 ));
defparam \instreth[20]~75 .lut_mask = 16'hA50A;
defparam \instreth[20]~75 .sum_lutc_input = "cin";

dffeas \instreth[20] (
	.clk(clock),
	.d(\instreth[20]~75_combout ),
	.asdata(\_T_244[20]~33_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[20]~q ),
	.prn(vcc));
defparam \instreth[20] .is_wysiwyg = "true";
defparam \instreth[20] .power_up = "low";

cyclone10lp_lcell_comb \instreth[21]~77 (
	.dataa(\instreth[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[20]~76 ),
	.combout(\instreth[21]~77_combout ),
	.cout(\instreth[21]~78 ));
defparam \instreth[21]~77 .lut_mask = 16'h5A5F;
defparam \instreth[21]~77 .sum_lutc_input = "cin";

dffeas \instreth[21] (
	.clk(clock),
	.d(\instreth[21]~77_combout ),
	.asdata(\_T_244[21]~35_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[21]~q ),
	.prn(vcc));
defparam \instreth[21] .is_wysiwyg = "true";
defparam \instreth[21] .power_up = "low";

cyclone10lp_lcell_comb \instreth[22]~79 (
	.dataa(\instreth[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[21]~78 ),
	.combout(\instreth[22]~79_combout ),
	.cout(\instreth[22]~80 ));
defparam \instreth[22]~79 .lut_mask = 16'hA50A;
defparam \instreth[22]~79 .sum_lutc_input = "cin";

dffeas \instreth[22] (
	.clk(clock),
	.d(\instreth[22]~79_combout ),
	.asdata(\_T_244[22]~37_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[22]~q ),
	.prn(vcc));
defparam \instreth[22] .is_wysiwyg = "true";
defparam \instreth[22] .power_up = "low";

cyclone10lp_lcell_comb \instreth[23]~81 (
	.dataa(\instreth[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[22]~80 ),
	.combout(\instreth[23]~81_combout ),
	.cout(\instreth[23]~82 ));
defparam \instreth[23]~81 .lut_mask = 16'h5A5F;
defparam \instreth[23]~81 .sum_lutc_input = "cin";

dffeas \instreth[23] (
	.clk(clock),
	.d(\instreth[23]~81_combout ),
	.asdata(\_T_244[23]~39_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[23]~q ),
	.prn(vcc));
defparam \instreth[23] .is_wysiwyg = "true";
defparam \instreth[23] .power_up = "low";

cyclone10lp_lcell_comb \instreth[24]~83 (
	.dataa(\instreth[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[23]~82 ),
	.combout(\instreth[24]~83_combout ),
	.cout(\instreth[24]~84 ));
defparam \instreth[24]~83 .lut_mask = 16'hA50A;
defparam \instreth[24]~83 .sum_lutc_input = "cin";

dffeas \instreth[24] (
	.clk(clock),
	.d(\instreth[24]~83_combout ),
	.asdata(\_T_244[24]~41_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[24]~q ),
	.prn(vcc));
defparam \instreth[24] .is_wysiwyg = "true";
defparam \instreth[24] .power_up = "low";

cyclone10lp_lcell_comb \instreth[25]~85 (
	.dataa(\instreth[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[24]~84 ),
	.combout(\instreth[25]~85_combout ),
	.cout(\instreth[25]~86 ));
defparam \instreth[25]~85 .lut_mask = 16'h5A5F;
defparam \instreth[25]~85 .sum_lutc_input = "cin";

dffeas \instreth[25] (
	.clk(clock),
	.d(\instreth[25]~85_combout ),
	.asdata(\_T_244[25]~43_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[25]~q ),
	.prn(vcc));
defparam \instreth[25] .is_wysiwyg = "true";
defparam \instreth[25] .power_up = "low";

cyclone10lp_lcell_comb \instreth[26]~87 (
	.dataa(\instreth[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[25]~86 ),
	.combout(\instreth[26]~87_combout ),
	.cout(\instreth[26]~88 ));
defparam \instreth[26]~87 .lut_mask = 16'hA50A;
defparam \instreth[26]~87 .sum_lutc_input = "cin";

dffeas \instreth[26] (
	.clk(clock),
	.d(\instreth[26]~87_combout ),
	.asdata(\_T_244[26]~45_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[26]~q ),
	.prn(vcc));
defparam \instreth[26] .is_wysiwyg = "true";
defparam \instreth[26] .power_up = "low";

cyclone10lp_lcell_comb \instreth[27]~89 (
	.dataa(\instreth[27]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[26]~88 ),
	.combout(\instreth[27]~89_combout ),
	.cout(\instreth[27]~90 ));
defparam \instreth[27]~89 .lut_mask = 16'h5A5F;
defparam \instreth[27]~89 .sum_lutc_input = "cin";

dffeas \instreth[27] (
	.clk(clock),
	.d(\instreth[27]~89_combout ),
	.asdata(\_T_244[27]~47_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[27]~q ),
	.prn(vcc));
defparam \instreth[27] .is_wysiwyg = "true";
defparam \instreth[27] .power_up = "low";

cyclone10lp_lcell_comb \instreth[28]~91 (
	.dataa(\instreth[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[27]~90 ),
	.combout(\instreth[28]~91_combout ),
	.cout(\instreth[28]~92 ));
defparam \instreth[28]~91 .lut_mask = 16'hA50A;
defparam \instreth[28]~91 .sum_lutc_input = "cin";

dffeas \instreth[28] (
	.clk(clock),
	.d(\instreth[28]~91_combout ),
	.asdata(\_T_244[28]~49_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[28]~q ),
	.prn(vcc));
defparam \instreth[28] .is_wysiwyg = "true";
defparam \instreth[28] .power_up = "low";

cyclone10lp_lcell_comb \io_out[28]~30 (
	.dataa(\io_out[1]~14_combout ),
	.datab(\instreth[28]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[28]~30_combout ),
	.cout());
defparam \io_out[28]~30 .lut_mask = 16'h8888;
defparam \io_out[28]~30 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \timeh[2]~40 (
	.dataa(\timeh[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[1]~37 ),
	.combout(\timeh[2]~40_combout ),
	.cout(\timeh[2]~41 ));
defparam \timeh[2]~40 .lut_mask = 16'hA50A;
defparam \timeh[2]~40 .sum_lutc_input = "cin";

dffeas \timeh[2] (
	.clk(clock),
	.d(\timeh[2]~40_combout ),
	.asdata(\_T_246[2]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[2]~q ),
	.prn(vcc));
defparam \timeh[2] .is_wysiwyg = "true";
defparam \timeh[2] .power_up = "low";

cyclone10lp_lcell_comb \timeh[3]~42 (
	.dataa(\timeh[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[2]~41 ),
	.combout(\timeh[3]~42_combout ),
	.cout(\timeh[3]~43 ));
defparam \timeh[3]~42 .lut_mask = 16'h5A5F;
defparam \timeh[3]~42 .sum_lutc_input = "cin";

dffeas \timeh[3] (
	.clk(clock),
	.d(\timeh[3]~42_combout ),
	.asdata(\_T_246[3]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[3]~q ),
	.prn(vcc));
defparam \timeh[3] .is_wysiwyg = "true";
defparam \timeh[3] .power_up = "low";

cyclone10lp_lcell_comb \timeh[4]~44 (
	.dataa(\timeh[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[3]~43 ),
	.combout(\timeh[4]~44_combout ),
	.cout(\timeh[4]~45 ));
defparam \timeh[4]~44 .lut_mask = 16'hA50A;
defparam \timeh[4]~44 .sum_lutc_input = "cin";

dffeas \timeh[4] (
	.clk(clock),
	.d(\timeh[4]~44_combout ),
	.asdata(\_T_244[4]~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[4]~q ),
	.prn(vcc));
defparam \timeh[4] .is_wysiwyg = "true";
defparam \timeh[4] .power_up = "low";

cyclone10lp_lcell_comb \timeh[5]~46 (
	.dataa(\timeh[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[4]~45 ),
	.combout(\timeh[5]~46_combout ),
	.cout(\timeh[5]~47 ));
defparam \timeh[5]~46 .lut_mask = 16'h5A5F;
defparam \timeh[5]~46 .sum_lutc_input = "cin";

dffeas \timeh[5] (
	.clk(clock),
	.d(\timeh[5]~46_combout ),
	.asdata(\_T_244[5]~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[5]~q ),
	.prn(vcc));
defparam \timeh[5] .is_wysiwyg = "true";
defparam \timeh[5] .power_up = "low";

cyclone10lp_lcell_comb \timeh[6]~48 (
	.dataa(\timeh[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[5]~47 ),
	.combout(\timeh[6]~48_combout ),
	.cout(\timeh[6]~49 ));
defparam \timeh[6]~48 .lut_mask = 16'hA50A;
defparam \timeh[6]~48 .sum_lutc_input = "cin";

dffeas \timeh[6] (
	.clk(clock),
	.d(\timeh[6]~48_combout ),
	.asdata(\_T_244[6]~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[6]~q ),
	.prn(vcc));
defparam \timeh[6] .is_wysiwyg = "true";
defparam \timeh[6] .power_up = "low";

cyclone10lp_lcell_comb \timeh[7]~50 (
	.dataa(\timeh[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[6]~49 ),
	.combout(\timeh[7]~50_combout ),
	.cout(\timeh[7]~51 ));
defparam \timeh[7]~50 .lut_mask = 16'h5A5F;
defparam \timeh[7]~50 .sum_lutc_input = "cin";

dffeas \timeh[7] (
	.clk(clock),
	.d(\timeh[7]~50_combout ),
	.asdata(\_T_244[7]~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[7]~q ),
	.prn(vcc));
defparam \timeh[7] .is_wysiwyg = "true";
defparam \timeh[7] .power_up = "low";

cyclone10lp_lcell_comb \timeh[8]~52 (
	.dataa(\timeh[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[7]~51 ),
	.combout(\timeh[8]~52_combout ),
	.cout(\timeh[8]~53 ));
defparam \timeh[8]~52 .lut_mask = 16'hA50A;
defparam \timeh[8]~52 .sum_lutc_input = "cin";

dffeas \timeh[8] (
	.clk(clock),
	.d(\timeh[8]~52_combout ),
	.asdata(\_T_244[8]~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[8]~q ),
	.prn(vcc));
defparam \timeh[8] .is_wysiwyg = "true";
defparam \timeh[8] .power_up = "low";

cyclone10lp_lcell_comb \timeh[9]~54 (
	.dataa(\timeh[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[8]~53 ),
	.combout(\timeh[9]~54_combout ),
	.cout(\timeh[9]~55 ));
defparam \timeh[9]~54 .lut_mask = 16'h5A5F;
defparam \timeh[9]~54 .sum_lutc_input = "cin";

dffeas \timeh[9] (
	.clk(clock),
	.d(\timeh[9]~54_combout ),
	.asdata(\_T_244[9]~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[9]~q ),
	.prn(vcc));
defparam \timeh[9] .is_wysiwyg = "true";
defparam \timeh[9] .power_up = "low";

cyclone10lp_lcell_comb \timeh[10]~56 (
	.dataa(\timeh[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[9]~55 ),
	.combout(\timeh[10]~56_combout ),
	.cout(\timeh[10]~57 ));
defparam \timeh[10]~56 .lut_mask = 16'hA50A;
defparam \timeh[10]~56 .sum_lutc_input = "cin";

dffeas \timeh[10] (
	.clk(clock),
	.d(\timeh[10]~56_combout ),
	.asdata(\_T_244[10]~13_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[10]~q ),
	.prn(vcc));
defparam \timeh[10] .is_wysiwyg = "true";
defparam \timeh[10] .power_up = "low";

cyclone10lp_lcell_comb \timeh[11]~58 (
	.dataa(\timeh[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[10]~57 ),
	.combout(\timeh[11]~58_combout ),
	.cout(\timeh[11]~59 ));
defparam \timeh[11]~58 .lut_mask = 16'h5A5F;
defparam \timeh[11]~58 .sum_lutc_input = "cin";

dffeas \timeh[11] (
	.clk(clock),
	.d(\timeh[11]~58_combout ),
	.asdata(\_T_244[11]~15_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[11]~q ),
	.prn(vcc));
defparam \timeh[11] .is_wysiwyg = "true";
defparam \timeh[11] .power_up = "low";

cyclone10lp_lcell_comb \timeh[12]~60 (
	.dataa(\timeh[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[11]~59 ),
	.combout(\timeh[12]~60_combout ),
	.cout(\timeh[12]~61 ));
defparam \timeh[12]~60 .lut_mask = 16'hA50A;
defparam \timeh[12]~60 .sum_lutc_input = "cin";

dffeas \timeh[12] (
	.clk(clock),
	.d(\timeh[12]~60_combout ),
	.asdata(\_T_244[12]~17_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[12]~q ),
	.prn(vcc));
defparam \timeh[12] .is_wysiwyg = "true";
defparam \timeh[12] .power_up = "low";

cyclone10lp_lcell_comb \timeh[13]~62 (
	.dataa(\timeh[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[12]~61 ),
	.combout(\timeh[13]~62_combout ),
	.cout(\timeh[13]~63 ));
defparam \timeh[13]~62 .lut_mask = 16'h5A5F;
defparam \timeh[13]~62 .sum_lutc_input = "cin";

dffeas \timeh[13] (
	.clk(clock),
	.d(\timeh[13]~62_combout ),
	.asdata(\_T_244[13]~19_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[13]~q ),
	.prn(vcc));
defparam \timeh[13] .is_wysiwyg = "true";
defparam \timeh[13] .power_up = "low";

cyclone10lp_lcell_comb \timeh[14]~64 (
	.dataa(\timeh[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[13]~63 ),
	.combout(\timeh[14]~64_combout ),
	.cout(\timeh[14]~65 ));
defparam \timeh[14]~64 .lut_mask = 16'hA50A;
defparam \timeh[14]~64 .sum_lutc_input = "cin";

dffeas \timeh[14] (
	.clk(clock),
	.d(\timeh[14]~64_combout ),
	.asdata(\_T_244[14]~21_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[14]~q ),
	.prn(vcc));
defparam \timeh[14] .is_wysiwyg = "true";
defparam \timeh[14] .power_up = "low";

cyclone10lp_lcell_comb \timeh[15]~66 (
	.dataa(\timeh[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[14]~65 ),
	.combout(\timeh[15]~66_combout ),
	.cout(\timeh[15]~67 ));
defparam \timeh[15]~66 .lut_mask = 16'h5A5F;
defparam \timeh[15]~66 .sum_lutc_input = "cin";

dffeas \timeh[15] (
	.clk(clock),
	.d(\timeh[15]~66_combout ),
	.asdata(\_T_244[15]~23_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[15]~q ),
	.prn(vcc));
defparam \timeh[15] .is_wysiwyg = "true";
defparam \timeh[15] .power_up = "low";

cyclone10lp_lcell_comb \timeh[16]~68 (
	.dataa(\timeh[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[15]~67 ),
	.combout(\timeh[16]~68_combout ),
	.cout(\timeh[16]~69 ));
defparam \timeh[16]~68 .lut_mask = 16'hA50A;
defparam \timeh[16]~68 .sum_lutc_input = "cin";

dffeas \timeh[16] (
	.clk(clock),
	.d(\timeh[16]~68_combout ),
	.asdata(\_T_244[16]~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[16]~q ),
	.prn(vcc));
defparam \timeh[16] .is_wysiwyg = "true";
defparam \timeh[16] .power_up = "low";

cyclone10lp_lcell_comb \timeh[17]~70 (
	.dataa(\timeh[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[16]~69 ),
	.combout(\timeh[17]~70_combout ),
	.cout(\timeh[17]~71 ));
defparam \timeh[17]~70 .lut_mask = 16'h5A5F;
defparam \timeh[17]~70 .sum_lutc_input = "cin";

dffeas \timeh[17] (
	.clk(clock),
	.d(\timeh[17]~70_combout ),
	.asdata(\_T_244[17]~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[17]~q ),
	.prn(vcc));
defparam \timeh[17] .is_wysiwyg = "true";
defparam \timeh[17] .power_up = "low";

cyclone10lp_lcell_comb \timeh[18]~72 (
	.dataa(\timeh[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[17]~71 ),
	.combout(\timeh[18]~72_combout ),
	.cout(\timeh[18]~73 ));
defparam \timeh[18]~72 .lut_mask = 16'hA50A;
defparam \timeh[18]~72 .sum_lutc_input = "cin";

dffeas \timeh[18] (
	.clk(clock),
	.d(\timeh[18]~72_combout ),
	.asdata(\_T_244[18]~29_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[18]~q ),
	.prn(vcc));
defparam \timeh[18] .is_wysiwyg = "true";
defparam \timeh[18] .power_up = "low";

cyclone10lp_lcell_comb \timeh[19]~74 (
	.dataa(\timeh[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[18]~73 ),
	.combout(\timeh[19]~74_combout ),
	.cout(\timeh[19]~75 ));
defparam \timeh[19]~74 .lut_mask = 16'h5A5F;
defparam \timeh[19]~74 .sum_lutc_input = "cin";

dffeas \timeh[19] (
	.clk(clock),
	.d(\timeh[19]~74_combout ),
	.asdata(\_T_244[19]~31_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[19]~q ),
	.prn(vcc));
defparam \timeh[19] .is_wysiwyg = "true";
defparam \timeh[19] .power_up = "low";

cyclone10lp_lcell_comb \timeh[20]~76 (
	.dataa(\timeh[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[19]~75 ),
	.combout(\timeh[20]~76_combout ),
	.cout(\timeh[20]~77 ));
defparam \timeh[20]~76 .lut_mask = 16'hA50A;
defparam \timeh[20]~76 .sum_lutc_input = "cin";

dffeas \timeh[20] (
	.clk(clock),
	.d(\timeh[20]~76_combout ),
	.asdata(\_T_244[20]~33_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[20]~q ),
	.prn(vcc));
defparam \timeh[20] .is_wysiwyg = "true";
defparam \timeh[20] .power_up = "low";

cyclone10lp_lcell_comb \timeh[21]~78 (
	.dataa(\timeh[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[20]~77 ),
	.combout(\timeh[21]~78_combout ),
	.cout(\timeh[21]~79 ));
defparam \timeh[21]~78 .lut_mask = 16'h5A5F;
defparam \timeh[21]~78 .sum_lutc_input = "cin";

dffeas \timeh[21] (
	.clk(clock),
	.d(\timeh[21]~78_combout ),
	.asdata(\_T_244[21]~35_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[21]~q ),
	.prn(vcc));
defparam \timeh[21] .is_wysiwyg = "true";
defparam \timeh[21] .power_up = "low";

cyclone10lp_lcell_comb \timeh[22]~80 (
	.dataa(\timeh[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[21]~79 ),
	.combout(\timeh[22]~80_combout ),
	.cout(\timeh[22]~81 ));
defparam \timeh[22]~80 .lut_mask = 16'hA50A;
defparam \timeh[22]~80 .sum_lutc_input = "cin";

dffeas \timeh[22] (
	.clk(clock),
	.d(\timeh[22]~80_combout ),
	.asdata(\_T_244[22]~37_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[22]~q ),
	.prn(vcc));
defparam \timeh[22] .is_wysiwyg = "true";
defparam \timeh[22] .power_up = "low";

cyclone10lp_lcell_comb \timeh[23]~82 (
	.dataa(\timeh[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[22]~81 ),
	.combout(\timeh[23]~82_combout ),
	.cout(\timeh[23]~83 ));
defparam \timeh[23]~82 .lut_mask = 16'h5A5F;
defparam \timeh[23]~82 .sum_lutc_input = "cin";

dffeas \timeh[23] (
	.clk(clock),
	.d(\timeh[23]~82_combout ),
	.asdata(\_T_244[23]~39_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[23]~q ),
	.prn(vcc));
defparam \timeh[23] .is_wysiwyg = "true";
defparam \timeh[23] .power_up = "low";

cyclone10lp_lcell_comb \timeh[24]~84 (
	.dataa(\timeh[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[23]~83 ),
	.combout(\timeh[24]~84_combout ),
	.cout(\timeh[24]~85 ));
defparam \timeh[24]~84 .lut_mask = 16'hA50A;
defparam \timeh[24]~84 .sum_lutc_input = "cin";

dffeas \timeh[24] (
	.clk(clock),
	.d(\timeh[24]~84_combout ),
	.asdata(\_T_244[24]~41_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[24]~q ),
	.prn(vcc));
defparam \timeh[24] .is_wysiwyg = "true";
defparam \timeh[24] .power_up = "low";

cyclone10lp_lcell_comb \timeh[25]~86 (
	.dataa(\timeh[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[24]~85 ),
	.combout(\timeh[25]~86_combout ),
	.cout(\timeh[25]~87 ));
defparam \timeh[25]~86 .lut_mask = 16'h5A5F;
defparam \timeh[25]~86 .sum_lutc_input = "cin";

dffeas \timeh[25] (
	.clk(clock),
	.d(\timeh[25]~86_combout ),
	.asdata(\_T_244[25]~43_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[25]~q ),
	.prn(vcc));
defparam \timeh[25] .is_wysiwyg = "true";
defparam \timeh[25] .power_up = "low";

cyclone10lp_lcell_comb \timeh[26]~88 (
	.dataa(\timeh[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[25]~87 ),
	.combout(\timeh[26]~88_combout ),
	.cout(\timeh[26]~89 ));
defparam \timeh[26]~88 .lut_mask = 16'hA50A;
defparam \timeh[26]~88 .sum_lutc_input = "cin";

dffeas \timeh[26] (
	.clk(clock),
	.d(\timeh[26]~88_combout ),
	.asdata(\_T_244[26]~45_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[26]~q ),
	.prn(vcc));
defparam \timeh[26] .is_wysiwyg = "true";
defparam \timeh[26] .power_up = "low";

cyclone10lp_lcell_comb \timeh[27]~90 (
	.dataa(\timeh[27]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[26]~89 ),
	.combout(\timeh[27]~90_combout ),
	.cout(\timeh[27]~91 ));
defparam \timeh[27]~90 .lut_mask = 16'h5A5F;
defparam \timeh[27]~90 .sum_lutc_input = "cin";

dffeas \timeh[27] (
	.clk(clock),
	.d(\timeh[27]~90_combout ),
	.asdata(\_T_244[27]~47_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[27]~q ),
	.prn(vcc));
defparam \timeh[27] .is_wysiwyg = "true";
defparam \timeh[27] .power_up = "low";

cyclone10lp_lcell_comb \timeh[28]~92 (
	.dataa(\timeh[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[27]~91 ),
	.combout(\timeh[28]~92_combout ),
	.cout(\timeh[28]~93 ));
defparam \timeh[28]~92 .lut_mask = 16'hA50A;
defparam \timeh[28]~92 .sum_lutc_input = "cin";

dffeas \timeh[28] (
	.clk(clock),
	.d(\timeh[28]~92_combout ),
	.asdata(\_T_244[28]~49_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[28]~q ),
	.prn(vcc));
defparam \timeh[28] .is_wysiwyg = "true";
defparam \timeh[28] .power_up = "low";

dffeas \mscratch[29] (
	.clk(clock),
	.d(\_T_244[29]~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[29]~q ),
	.prn(vcc));
defparam \mscratch[29] .is_wysiwyg = "true";
defparam \mscratch[29] .power_up = "low";

cyclone10lp_lcell_comb \io_out[29]~32 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[29]~q ),
	.datad(\mscratch[29]~q ),
	.cin(gnd),
	.combout(\io_out[29]~32_combout ),
	.cout());
defparam \io_out[29]~32 .lut_mask = 16'hEAC0;
defparam \io_out[29]~32 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[29]~33 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_29),
	.datad(\time_[29]~q ),
	.cin(gnd),
	.combout(\io_out[29]~33_combout ),
	.cout());
defparam \io_out[29]~33 .lut_mask = 16'hEAC0;
defparam \io_out[29]~33 .sum_lutc_input = "datac";

dffeas \mbadaddr[29] (
	.clk(clock),
	.d(\_T_244[29]~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[29]~q ),
	.prn(vcc));
defparam \mbadaddr[29] .is_wysiwyg = "true";
defparam \mbadaddr[29] .power_up = "low";

cyclone10lp_lcell_comb \io_out[29]~34 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[29]~q ),
	.datad(\mbadaddr[29]~q ),
	.cin(gnd),
	.combout(\io_out[29]~34_combout ),
	.cout());
defparam \io_out[29]~34 .lut_mask = 16'hEAC0;
defparam \io_out[29]~34 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cycleh[29]~92 (
	.dataa(\cycleh[29]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[28]~91 ),
	.combout(\cycleh[29]~92_combout ),
	.cout(\cycleh[29]~93 ));
defparam \cycleh[29]~92 .lut_mask = 16'h5A5F;
defparam \cycleh[29]~92 .sum_lutc_input = "cin";

dffeas \cycleh[29] (
	.clk(clock),
	.d(\cycleh[29]~92_combout ),
	.asdata(\_T_244[29]~51_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[29]~q ),
	.prn(vcc));
defparam \cycleh[29] .is_wysiwyg = "true";
defparam \cycleh[29] .power_up = "low";

cyclone10lp_lcell_comb \io_out[29]~35 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_29),
	.datad(\cycleh[29]~q ),
	.cin(gnd),
	.combout(\io_out[29]~35_combout ),
	.cout());
defparam \io_out[29]~35 .lut_mask = 16'hEAC0;
defparam \io_out[29]~35 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \instreth[29]~93 (
	.dataa(\instreth[29]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[28]~92 ),
	.combout(\instreth[29]~93_combout ),
	.cout(\instreth[29]~94 ));
defparam \instreth[29]~93 .lut_mask = 16'h5A5F;
defparam \instreth[29]~93 .sum_lutc_input = "cin";

dffeas \instreth[29] (
	.clk(clock),
	.d(\instreth[29]~93_combout ),
	.asdata(\_T_244[29]~51_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[29]~q ),
	.prn(vcc));
defparam \instreth[29] .is_wysiwyg = "true";
defparam \instreth[29] .power_up = "low";

cyclone10lp_lcell_comb \timeh[29]~94 (
	.dataa(\timeh[29]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[28]~93 ),
	.combout(\timeh[29]~94_combout ),
	.cout(\timeh[29]~95 ));
defparam \timeh[29]~94 .lut_mask = 16'h5A5F;
defparam \timeh[29]~94 .sum_lutc_input = "cin";

dffeas \timeh[29] (
	.clk(clock),
	.d(\timeh[29]~94_combout ),
	.asdata(\_T_244[29]~51_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[29]~q ),
	.prn(vcc));
defparam \timeh[29] .is_wysiwyg = "true";
defparam \timeh[29] .power_up = "low";

dffeas \mscratch[30] (
	.clk(clock),
	.d(\_T_244[30]~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[30]~q ),
	.prn(vcc));
defparam \mscratch[30] .is_wysiwyg = "true";
defparam \mscratch[30] .power_up = "low";

cyclone10lp_lcell_comb \io_out[30]~39 (
	.dataa(\Equal25~5_combout ),
	.datab(\Equal25~3_combout ),
	.datac(\mscratch[30]~q ),
	.datad(\Equal19~2_combout ),
	.cin(gnd),
	.combout(\io_out[30]~39_combout ),
	.cout());
defparam \io_out[30]~39 .lut_mask = 16'hEAC0;
defparam \io_out[30]~39 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[30]~40 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_30),
	.datad(\time_[30]~q ),
	.cin(gnd),
	.combout(\io_out[30]~40_combout ),
	.cout());
defparam \io_out[30]~40 .lut_mask = 16'hEAC0;
defparam \io_out[30]~40 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[30]~41 (
	.dataa(\io_out[30]~39_combout ),
	.datab(\io_out[30]~40_combout ),
	.datac(\io_out[1]~6_combout ),
	.datad(\cycle[30]~q ),
	.cin(gnd),
	.combout(\io_out[30]~41_combout ),
	.cout());
defparam \io_out[30]~41 .lut_mask = 16'hFEEE;
defparam \io_out[30]~41 .sum_lutc_input = "datac";

dffeas \mbadaddr[30] (
	.clk(clock),
	.d(\_T_244[30]~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[30]~q ),
	.prn(vcc));
defparam \mbadaddr[30] .is_wysiwyg = "true";
defparam \mbadaddr[30] .power_up = "low";

cyclone10lp_lcell_comb \io_out[30]~42 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[30]~q ),
	.datad(\mbadaddr[30]~q ),
	.cin(gnd),
	.combout(\io_out[30]~42_combout ),
	.cout());
defparam \io_out[30]~42 .lut_mask = 16'hEAC0;
defparam \io_out[30]~42 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cycleh[30]~94 (
	.dataa(\cycleh[30]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\cycleh[29]~93 ),
	.combout(\cycleh[30]~94_combout ),
	.cout(\cycleh[30]~95 ));
defparam \cycleh[30]~94 .lut_mask = 16'hA50A;
defparam \cycleh[30]~94 .sum_lutc_input = "cin";

dffeas \cycleh[30] (
	.clk(clock),
	.d(\cycleh[30]~94_combout ),
	.asdata(\_T_244[30]~53_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[30]~q ),
	.prn(vcc));
defparam \cycleh[30] .is_wysiwyg = "true";
defparam \cycleh[30] .power_up = "low";

cyclone10lp_lcell_comb \io_out[30]~43 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_30),
	.datad(\cycleh[30]~q ),
	.cin(gnd),
	.combout(\io_out[30]~43_combout ),
	.cout());
defparam \io_out[30]~43 .lut_mask = 16'hEAC0;
defparam \io_out[30]~43 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \instreth[30]~95 (
	.dataa(\instreth[30]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\instreth[29]~94 ),
	.combout(\instreth[30]~95_combout ),
	.cout(\instreth[30]~96 ));
defparam \instreth[30]~95 .lut_mask = 16'hA50A;
defparam \instreth[30]~95 .sum_lutc_input = "cin";

dffeas \instreth[30] (
	.clk(clock),
	.d(\instreth[30]~95_combout ),
	.asdata(\_T_244[30]~53_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[30]~q ),
	.prn(vcc));
defparam \instreth[30] .is_wysiwyg = "true";
defparam \instreth[30] .power_up = "low";

cyclone10lp_lcell_comb \timeh[30]~96 (
	.dataa(\timeh[30]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\timeh[29]~95 ),
	.combout(\timeh[30]~96_combout ),
	.cout(\timeh[30]~97 ));
defparam \timeh[30]~96 .lut_mask = 16'hA50A;
defparam \timeh[30]~96 .sum_lutc_input = "cin";

dffeas \timeh[30] (
	.clk(clock),
	.d(\timeh[30]~96_combout ),
	.asdata(\_T_244[30]~53_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[30]~q ),
	.prn(vcc));
defparam \timeh[30] .is_wysiwyg = "true";
defparam \timeh[30] .power_up = "low";

cyclone10lp_lcell_comb \io_out[30]~44 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[30]~q ),
	.datad(\timeh[30]~q ),
	.cin(gnd),
	.combout(\io_out[30]~44_combout ),
	.cout());
defparam \io_out[30]~44 .lut_mask = 16'hEAC0;
defparam \io_out[30]~44 .sum_lutc_input = "datac";

dffeas \mscratch[31] (
	.clk(clock),
	.d(\_T_246[31]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[31]~q ),
	.prn(vcc));
defparam \mscratch[31] .is_wysiwyg = "true";
defparam \mscratch[31] .power_up = "low";

cyclone10lp_lcell_comb \io_out[31]~46 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[31]~q ),
	.datad(\mscratch[31]~q ),
	.cin(gnd),
	.combout(\io_out[31]~46_combout ),
	.cout());
defparam \io_out[31]~46 .lut_mask = 16'hEAC0;
defparam \io_out[31]~46 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[31]~47 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_31),
	.datad(\time_[31]~q ),
	.cin(gnd),
	.combout(\io_out[31]~47_combout ),
	.cout());
defparam \io_out[31]~47 .lut_mask = 16'hEAC0;
defparam \io_out[31]~47 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mcause[31]~13 (
	.dataa(io_expt1),
	.datab(\_T_246[31]~10_combout ),
	.datac(gnd),
	.datad(isEcall),
	.cin(gnd),
	.combout(\mcause[31]~13_combout ),
	.cout());
defparam \mcause[31]~13 .lut_mask = 16'h0088;
defparam \mcause[31]~13 .sum_lutc_input = "datac";

dffeas \mcause[31] (
	.clk(clock),
	.d(\mcause[31]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mcause[0]~11_combout ),
	.q(\mcause[31]~q ),
	.prn(vcc));
defparam \mcause[31] .is_wysiwyg = "true";
defparam \mcause[31] .power_up = "low";

cyclone10lp_lcell_comb \io_out[31]~48 (
	.dataa(\Equal27~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[31]~q ),
	.datad(\mcause[31]~q ),
	.cin(gnd),
	.combout(\io_out[31]~48_combout ),
	.cout());
defparam \io_out[31]~48 .lut_mask = 16'hEAC0;
defparam \io_out[31]~48 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \cycleh[31]~96 (
	.dataa(\cycleh[31]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\cycleh[30]~95 ),
	.combout(\cycleh[31]~96_combout ),
	.cout());
defparam \cycleh[31]~96 .lut_mask = 16'h5A5A;
defparam \cycleh[31]~96 .sum_lutc_input = "cin";

dffeas \cycleh[31] (
	.clk(clock),
	.d(\cycleh[31]~96_combout ),
	.asdata(\_T_246[31]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\cycleh~36_combout ),
	.ena(\cycleh[23]~37_combout ),
	.q(\cycleh[31]~q ),
	.prn(vcc));
defparam \cycleh[31] .is_wysiwyg = "true";
defparam \cycleh[31] .power_up = "low";

dffeas \mbadaddr[31] (
	.clk(clock),
	.d(\_T_246[31]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[31]~q ),
	.prn(vcc));
defparam \mbadaddr[31] .is_wysiwyg = "true";
defparam \mbadaddr[31] .power_up = "low";

cyclone10lp_lcell_comb \io_out[31]~49 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~10_combout ),
	.datac(\cycleh[31]~q ),
	.datad(\mbadaddr[31]~q ),
	.cin(gnd),
	.combout(\io_out[31]~49_combout ),
	.cout());
defparam \io_out[31]~49 .lut_mask = 16'hEAC0;
defparam \io_out[31]~49 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[31]~50 (
	.dataa(\io_out[31]~46_combout ),
	.datab(\io_out[31]~47_combout ),
	.datac(\io_out[31]~48_combout ),
	.datad(\io_out[31]~49_combout ),
	.cin(gnd),
	.combout(\io_out[31]~50_combout ),
	.cout());
defparam \io_out[31]~50 .lut_mask = 16'hFFFE;
defparam \io_out[31]~50 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \timeh[31]~98 (
	.dataa(\timeh[31]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\timeh[30]~97 ),
	.combout(\timeh[31]~98_combout ),
	.cout());
defparam \timeh[31]~98 .lut_mask = 16'h5A5A;
defparam \timeh[31]~98 .sum_lutc_input = "cin";

dffeas \timeh[31] (
	.clk(clock),
	.d(\timeh[31]~98_combout ),
	.asdata(\_T_246[31]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\timeh~38_combout ),
	.ena(\timeh[31]~39_combout ),
	.q(\timeh[31]~q ),
	.prn(vcc));
defparam \timeh[31] .is_wysiwyg = "true";
defparam \timeh[31] .power_up = "low";

cyclone10lp_lcell_comb \io_out[31]~51 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_31),
	.datad(\timeh[31]~q ),
	.cin(gnd),
	.combout(\io_out[31]~51_combout ),
	.cout());
defparam \io_out[31]~51 .lut_mask = 16'hEAC0;
defparam \io_out[31]~51 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \instreth[31]~97 (
	.dataa(\instreth[31]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\instreth[30]~96 ),
	.combout(\instreth[31]~97_combout ),
	.cout());
defparam \instreth[31]~97 .lut_mask = 16'h5A5A;
defparam \instreth[31]~97 .sum_lutc_input = "cin";

dffeas \instreth[31] (
	.clk(clock),
	.d(\instreth[31]~97_combout ),
	.asdata(\_T_246[31]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(\instreth~37_combout ),
	.ena(\instreth[3]~38_combout ),
	.q(\instreth[31]~q ),
	.prn(vcc));
defparam \instreth[31] .is_wysiwyg = "true";
defparam \instreth[31] .power_up = "low";

cyclone10lp_lcell_comb \Equal16~2 (
	.dataa(Equal62),
	.datab(ex_csr_addr_10),
	.datac(\Equal16~0_combout ),
	.datad(\Equal16~1_combout ),
	.cin(gnd),
	.combout(\Equal16~2_combout ),
	.cout());
defparam \Equal16~2 .lut_mask = 16'h8000;
defparam \Equal16~2 .sum_lutc_input = "datac";

dffeas \mscratch[8] (
	.clk(clock),
	.d(\_T_244[8]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[8]~q ),
	.prn(vcc));
defparam \mscratch[8] .is_wysiwyg = "true";
defparam \mscratch[8] .power_up = "low";

cyclone10lp_lcell_comb \io_out[8]~53 (
	.dataa(\Equal16~2_combout ),
	.datab(\Equal25~3_combout ),
	.datac(\mscratch[8]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[8]~53_combout ),
	.cout());
defparam \io_out[8]~53 .lut_mask = 16'hEAEA;
defparam \io_out[8]~53 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[8]~54 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_8),
	.datad(\time_[8]~q ),
	.cin(gnd),
	.combout(\io_out[8]~54_combout ),
	.cout());
defparam \io_out[8]~54 .lut_mask = 16'hEAC0;
defparam \io_out[8]~54 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[8]~55 (
	.dataa(\io_out[8]~53_combout ),
	.datab(\io_out[8]~54_combout ),
	.datac(\io_out[1]~6_combout ),
	.datad(\cycle[8]~q ),
	.cin(gnd),
	.combout(\io_out[8]~55_combout ),
	.cout());
defparam \io_out[8]~55 .lut_mask = 16'hFEEE;
defparam \io_out[8]~55 .sum_lutc_input = "datac";

dffeas \mbadaddr[8] (
	.clk(clock),
	.d(\_T_244[8]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[8]~q ),
	.prn(vcc));
defparam \mbadaddr[8] .is_wysiwyg = "true";
defparam \mbadaddr[8] .power_up = "low";

cyclone10lp_lcell_comb \io_out[8]~56 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[8]~q ),
	.datad(\mbadaddr[8]~q ),
	.cin(gnd),
	.combout(\io_out[8]~56_combout ),
	.cout());
defparam \io_out[8]~56 .lut_mask = 16'hEAC0;
defparam \io_out[8]~56 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[8]~57 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_8),
	.datad(\cycleh[8]~q ),
	.cin(gnd),
	.combout(\io_out[8]~57_combout ),
	.cout());
defparam \io_out[8]~57 .lut_mask = 16'hEAC0;
defparam \io_out[8]~57 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[8]~58 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[8]~q ),
	.datad(\timeh[8]~q ),
	.cin(gnd),
	.combout(\io_out[8]~58_combout ),
	.cout());
defparam \io_out[8]~58 .lut_mask = 16'hEAC0;
defparam \io_out[8]~58 .sum_lutc_input = "datac";

dffeas \mscratch[9] (
	.clk(clock),
	.d(\_T_244[9]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[9]~q ),
	.prn(vcc));
defparam \mscratch[9] .is_wysiwyg = "true";
defparam \mscratch[9] .power_up = "low";

cyclone10lp_lcell_comb \io_out[9]~60 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[9]~q ),
	.datad(\mscratch[9]~q ),
	.cin(gnd),
	.combout(\io_out[9]~60_combout ),
	.cout());
defparam \io_out[9]~60 .lut_mask = 16'hEAC0;
defparam \io_out[9]~60 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[9]~61 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_9),
	.datad(\time_[9]~q ),
	.cin(gnd),
	.combout(\io_out[9]~61_combout ),
	.cout());
defparam \io_out[9]~61 .lut_mask = 16'hEAC0;
defparam \io_out[9]~61 .sum_lutc_input = "datac";

dffeas \mbadaddr[9] (
	.clk(clock),
	.d(\_T_244[9]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[9]~q ),
	.prn(vcc));
defparam \mbadaddr[9] .is_wysiwyg = "true";
defparam \mbadaddr[9] .power_up = "low";

cyclone10lp_lcell_comb \io_out[9]~62 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[9]~q ),
	.datad(\mbadaddr[9]~q ),
	.cin(gnd),
	.combout(\io_out[9]~62_combout ),
	.cout());
defparam \io_out[9]~62 .lut_mask = 16'hEAC0;
defparam \io_out[9]~62 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[9]~63 (
	.dataa(\Equal19~2_combout ),
	.datab(\Equal19~4_combout ),
	.datac(mtvec_9),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[9]~63_combout ),
	.cout());
defparam \io_out[9]~63 .lut_mask = 16'h8080;
defparam \io_out[9]~63 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[9]~64 (
	.dataa(\io_out[9]~62_combout ),
	.datab(\io_out[9]~63_combout ),
	.datac(\io_out[1]~10_combout ),
	.datad(\cycleh[9]~q ),
	.cin(gnd),
	.combout(\io_out[9]~64_combout ),
	.cout());
defparam \io_out[9]~64 .lut_mask = 16'hFEEE;
defparam \io_out[9]~64 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[9]~65 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[9]~q ),
	.datad(\timeh[9]~q ),
	.cin(gnd),
	.combout(\io_out[9]~65_combout ),
	.cout());
defparam \io_out[9]~65 .lut_mask = 16'hEAC0;
defparam \io_out[9]~65 .sum_lutc_input = "datac";

dffeas \mscratch[10] (
	.clk(clock),
	.d(\_T_244[10]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[10]~q ),
	.prn(vcc));
defparam \mscratch[10] .is_wysiwyg = "true";
defparam \mscratch[10] .power_up = "low";

cyclone10lp_lcell_comb \io_out[10]~67 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[10]~q ),
	.datad(\mscratch[10]~q ),
	.cin(gnd),
	.combout(\io_out[10]~67_combout ),
	.cout());
defparam \io_out[10]~67 .lut_mask = 16'hEAC0;
defparam \io_out[10]~67 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \Equal25~4 (
	.dataa(ex_csr_addr_6),
	.datab(\Equal25~2_combout ),
	.datac(\Equal16~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal25~4_combout ),
	.cout());
defparam \Equal25~4 .lut_mask = 16'h8080;
defparam \Equal25~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[10]~238 (
	.dataa(ex_csr_addr_0),
	.datab(ex_csr_addr_1),
	.datac(\Equal25~4_combout ),
	.datad(mepc_10),
	.cin(gnd),
	.combout(\io_out[10]~238_combout ),
	.cout());
defparam \io_out[10]~238 .lut_mask = 16'h2000;
defparam \io_out[10]~238 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[10]~68 (
	.dataa(\io_out[10]~67_combout ),
	.datab(\io_out[10]~238_combout ),
	.datac(\io_out[1]~4_combout ),
	.datad(\time_[10]~q ),
	.cin(gnd),
	.combout(\io_out[10]~68_combout ),
	.cout());
defparam \io_out[10]~68 .lut_mask = 16'hFEEE;
defparam \io_out[10]~68 .sum_lutc_input = "datac";

dffeas \mbadaddr[10] (
	.clk(clock),
	.d(\_T_244[10]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[10]~q ),
	.prn(vcc));
defparam \mbadaddr[10] .is_wysiwyg = "true";
defparam \mbadaddr[10] .power_up = "low";

cyclone10lp_lcell_comb \io_out[10]~69 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[10]~q ),
	.datad(\mbadaddr[10]~q ),
	.cin(gnd),
	.combout(\io_out[10]~69_combout ),
	.cout());
defparam \io_out[10]~69 .lut_mask = 16'hEAC0;
defparam \io_out[10]~69 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[10]~70 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_10),
	.datad(\cycleh[10]~q ),
	.cin(gnd),
	.combout(\io_out[10]~70_combout ),
	.cout());
defparam \io_out[10]~70 .lut_mask = 16'hEAC0;
defparam \io_out[10]~70 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[10]~71 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[10]~q ),
	.datad(\timeh[10]~q ),
	.cin(gnd),
	.combout(\io_out[10]~71_combout ),
	.cout());
defparam \io_out[10]~71 .lut_mask = 16'hEAC0;
defparam \io_out[10]~71 .sum_lutc_input = "datac";

dffeas \mscratch[11] (
	.clk(clock),
	.d(\_T_244[11]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[11]~q ),
	.prn(vcc));
defparam \mscratch[11] .is_wysiwyg = "true";
defparam \mscratch[11] .power_up = "low";

cyclone10lp_lcell_comb \io_out[11]~73 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~4_combout ),
	.datac(\time_[11]~q ),
	.datad(\mscratch[11]~q ),
	.cin(gnd),
	.combout(\io_out[11]~73_combout ),
	.cout());
defparam \io_out[11]~73 .lut_mask = 16'hEAC0;
defparam \io_out[11]~73 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[11]~74 (
	.dataa(\Equal26~0_combout ),
	.datab(\io_out[1]~12_combout ),
	.datac(\timeh[11]~q ),
	.datad(mepc_11),
	.cin(gnd),
	.combout(\io_out[11]~74_combout ),
	.cout());
defparam \io_out[11]~74 .lut_mask = 16'hEAC0;
defparam \io_out[11]~74 .sum_lutc_input = "datac";

dffeas \mbadaddr[11] (
	.clk(clock),
	.d(\_T_244[11]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[11]~q ),
	.prn(vcc));
defparam \mbadaddr[11] .is_wysiwyg = "true";
defparam \mbadaddr[11] .power_up = "low";

cyclone10lp_lcell_comb \io_out[11]~75 (
	.dataa(\io_out[1]~6_combout ),
	.datab(\Equal28~0_combout ),
	.datac(\mbadaddr[11]~q ),
	.datad(\cycle[11]~q ),
	.cin(gnd),
	.combout(\io_out[11]~75_combout ),
	.cout());
defparam \io_out[11]~75 .lut_mask = 16'hEAC0;
defparam \io_out[11]~75 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MTIE~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(gnd),
	.datac(\instreth~32_combout ),
	.datad(\Equal21~2_combout ),
	.cin(gnd),
	.combout(\MTIE~0_combout ),
	.cout());
defparam \MTIE~0 .lut_mask = 16'hF555;
defparam \MTIE~0 .sum_lutc_input = "datac";

dffeas MEIE(
	.clk(clock),
	.d(\mtvec~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MTIE~0_combout ),
	.q(\MEIE~q ),
	.prn(vcc));
defparam MEIE.is_wysiwyg = "true";
defparam MEIE.power_up = "low";

cyclone10lp_lcell_comb \io_out[11]~76 (
	.dataa(\Equal19~3_combout ),
	.datab(\Equal21~2_combout ),
	.datac(\MEIE~q ),
	.datad(mtvec_11),
	.cin(gnd),
	.combout(\io_out[11]~76_combout ),
	.cout());
defparam \io_out[11]~76 .lut_mask = 16'hEAC0;
defparam \io_out[11]~76 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[11]~77 (
	.dataa(\io_out[11]~75_combout ),
	.datab(\io_out[11]~76_combout ),
	.datac(\io_out[1]~8_combout ),
	.datad(\instret[11]~q ),
	.cin(gnd),
	.combout(\io_out[11]~77_combout ),
	.cout());
defparam \io_out[11]~77 .lut_mask = 16'hFEEE;
defparam \io_out[11]~77 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[11]~78 (
	.dataa(\io_out[1]~14_combout ),
	.datab(\io_out[1]~10_combout ),
	.datac(\cycleh[11]~q ),
	.datad(\instreth[11]~q ),
	.cin(gnd),
	.combout(\io_out[11]~78_combout ),
	.cout());
defparam \io_out[11]~78 .lut_mask = 16'hEAC0;
defparam \io_out[11]~78 .sum_lutc_input = "datac";

dffeas \mscratch[12] (
	.clk(clock),
	.d(\_T_244[12]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[12]~q ),
	.prn(vcc));
defparam \mscratch[12] .is_wysiwyg = "true";
defparam \mscratch[12] .power_up = "low";

cyclone10lp_lcell_comb \io_out[12]~80 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[12]~q ),
	.datad(\mscratch[12]~q ),
	.cin(gnd),
	.combout(\io_out[12]~80_combout ),
	.cout());
defparam \io_out[12]~80 .lut_mask = 16'hEAC0;
defparam \io_out[12]~80 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[12]~81 (
	.dataa(ex_csr_addr_6),
	.datab(\Equal25~5_combout ),
	.datac(\Equal4~0_combout ),
	.datad(mepc_12),
	.cin(gnd),
	.combout(\io_out[12]~81_combout ),
	.cout());
defparam \io_out[12]~81 .lut_mask = 16'h8000;
defparam \io_out[12]~81 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[12]~82 (
	.dataa(\io_out[12]~80_combout ),
	.datab(\io_out[12]~81_combout ),
	.datac(\io_out[1]~4_combout ),
	.datad(\time_[12]~q ),
	.cin(gnd),
	.combout(\io_out[12]~82_combout ),
	.cout());
defparam \io_out[12]~82 .lut_mask = 16'hFEEE;
defparam \io_out[12]~82 .sum_lutc_input = "datac";

dffeas \mbadaddr[12] (
	.clk(clock),
	.d(\_T_244[12]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[12]~q ),
	.prn(vcc));
defparam \mbadaddr[12] .is_wysiwyg = "true";
defparam \mbadaddr[12] .power_up = "low";

cyclone10lp_lcell_comb \io_out[12]~83 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[12]~q ),
	.datad(\mbadaddr[12]~q ),
	.cin(gnd),
	.combout(\io_out[12]~83_combout ),
	.cout());
defparam \io_out[12]~83 .lut_mask = 16'hEAC0;
defparam \io_out[12]~83 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[12]~84 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_12),
	.datad(\cycleh[12]~q ),
	.cin(gnd),
	.combout(\io_out[12]~84_combout ),
	.cout());
defparam \io_out[12]~84 .lut_mask = 16'hEAC0;
defparam \io_out[12]~84 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[12]~85 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[12]~q ),
	.datad(\timeh[12]~q ),
	.cin(gnd),
	.combout(\io_out[12]~85_combout ),
	.cout());
defparam \io_out[12]~85 .lut_mask = 16'hEAC0;
defparam \io_out[12]~85 .sum_lutc_input = "datac";

dffeas \mscratch[13] (
	.clk(clock),
	.d(\_T_244[13]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[13]~q ),
	.prn(vcc));
defparam \mscratch[13] .is_wysiwyg = "true";
defparam \mscratch[13] .power_up = "low";

cyclone10lp_lcell_comb \io_out[13]~87 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[13]~q ),
	.datad(\mscratch[13]~q ),
	.cin(gnd),
	.combout(\io_out[13]~87_combout ),
	.cout());
defparam \io_out[13]~87 .lut_mask = 16'hEAC0;
defparam \io_out[13]~87 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[13]~88 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_13),
	.datad(\time_[13]~q ),
	.cin(gnd),
	.combout(\io_out[13]~88_combout ),
	.cout());
defparam \io_out[13]~88 .lut_mask = 16'hEAC0;
defparam \io_out[13]~88 .sum_lutc_input = "datac";

dffeas \mbadaddr[13] (
	.clk(clock),
	.d(\_T_244[13]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[13]~q ),
	.prn(vcc));
defparam \mbadaddr[13] .is_wysiwyg = "true";
defparam \mbadaddr[13] .power_up = "low";

cyclone10lp_lcell_comb \io_out[13]~89 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[13]~q ),
	.datad(\mbadaddr[13]~q ),
	.cin(gnd),
	.combout(\io_out[13]~89_combout ),
	.cout());
defparam \io_out[13]~89 .lut_mask = 16'hEAC0;
defparam \io_out[13]~89 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[13]~90 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_13),
	.datad(\cycleh[13]~q ),
	.cin(gnd),
	.combout(\io_out[13]~90_combout ),
	.cout());
defparam \io_out[13]~90 .lut_mask = 16'hEAC0;
defparam \io_out[13]~90 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[13]~91 (
	.dataa(\io_out[13]~87_combout ),
	.datab(\io_out[13]~88_combout ),
	.datac(\io_out[13]~89_combout ),
	.datad(\io_out[13]~90_combout ),
	.cin(gnd),
	.combout(\io_out[13]~91_combout ),
	.cout());
defparam \io_out[13]~91 .lut_mask = 16'hFFFE;
defparam \io_out[13]~91 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[13]~92 (
	.dataa(\io_out[1]~14_combout ),
	.datab(\instreth[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[13]~92_combout ),
	.cout());
defparam \io_out[13]~92 .lut_mask = 16'h8888;
defparam \io_out[13]~92 .sum_lutc_input = "datac";

dffeas \mscratch[14] (
	.clk(clock),
	.d(\_T_244[14]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[14]~q ),
	.prn(vcc));
defparam \mscratch[14] .is_wysiwyg = "true";
defparam \mscratch[14] .power_up = "low";

cyclone10lp_lcell_comb \io_out[14]~94 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[14]~q ),
	.datad(\mscratch[14]~q ),
	.cin(gnd),
	.combout(\io_out[14]~94_combout ),
	.cout());
defparam \io_out[14]~94 .lut_mask = 16'hEAC0;
defparam \io_out[14]~94 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[14]~95 (
	.dataa(ex_csr_addr_0),
	.datab(\Equal25~4_combout ),
	.datac(mepc_14),
	.datad(ex_csr_addr_1),
	.cin(gnd),
	.combout(\io_out[14]~95_combout ),
	.cout());
defparam \io_out[14]~95 .lut_mask = 16'h0080;
defparam \io_out[14]~95 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[14]~96 (
	.dataa(\io_out[14]~94_combout ),
	.datab(\io_out[14]~95_combout ),
	.datac(\io_out[1]~4_combout ),
	.datad(\time_[14]~q ),
	.cin(gnd),
	.combout(\io_out[14]~96_combout ),
	.cout());
defparam \io_out[14]~96 .lut_mask = 16'hFEEE;
defparam \io_out[14]~96 .sum_lutc_input = "datac";

dffeas \mbadaddr[14] (
	.clk(clock),
	.d(\_T_244[14]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[14]~q ),
	.prn(vcc));
defparam \mbadaddr[14] .is_wysiwyg = "true";
defparam \mbadaddr[14] .power_up = "low";

cyclone10lp_lcell_comb \io_out[14]~97 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[14]~q ),
	.datad(\mbadaddr[14]~q ),
	.cin(gnd),
	.combout(\io_out[14]~97_combout ),
	.cout());
defparam \io_out[14]~97 .lut_mask = 16'hEAC0;
defparam \io_out[14]~97 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[14]~98 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_14),
	.datad(\cycleh[14]~q ),
	.cin(gnd),
	.combout(\io_out[14]~98_combout ),
	.cout());
defparam \io_out[14]~98 .lut_mask = 16'hEAC0;
defparam \io_out[14]~98 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[14]~99 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[14]~q ),
	.datad(\timeh[14]~q ),
	.cin(gnd),
	.combout(\io_out[14]~99_combout ),
	.cout());
defparam \io_out[14]~99 .lut_mask = 16'hEAC0;
defparam \io_out[14]~99 .sum_lutc_input = "datac";

dffeas \mscratch[15] (
	.clk(clock),
	.d(\_T_244[15]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[15]~q ),
	.prn(vcc));
defparam \mscratch[15] .is_wysiwyg = "true";
defparam \mscratch[15] .power_up = "low";

cyclone10lp_lcell_comb \io_out[15]~101 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[15]~q ),
	.datad(\mscratch[15]~q ),
	.cin(gnd),
	.combout(\io_out[15]~101_combout ),
	.cout());
defparam \io_out[15]~101 .lut_mask = 16'hEAC0;
defparam \io_out[15]~101 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[15]~102 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_15),
	.datad(\time_[15]~q ),
	.cin(gnd),
	.combout(\io_out[15]~102_combout ),
	.cout());
defparam \io_out[15]~102 .lut_mask = 16'hEAC0;
defparam \io_out[15]~102 .sum_lutc_input = "datac";

dffeas \mbadaddr[15] (
	.clk(clock),
	.d(\_T_244[15]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[15]~q ),
	.prn(vcc));
defparam \mbadaddr[15] .is_wysiwyg = "true";
defparam \mbadaddr[15] .power_up = "low";

cyclone10lp_lcell_comb \io_out[15]~103 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[15]~q ),
	.datad(\mbadaddr[15]~q ),
	.cin(gnd),
	.combout(\io_out[15]~103_combout ),
	.cout());
defparam \io_out[15]~103 .lut_mask = 16'hEAC0;
defparam \io_out[15]~103 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[15]~104 (
	.dataa(\Equal19~3_combout ),
	.datab(mtvec_15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[15]~104_combout ),
	.cout());
defparam \io_out[15]~104 .lut_mask = 16'h8888;
defparam \io_out[15]~104 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[15]~105 (
	.dataa(\io_out[15]~103_combout ),
	.datab(\io_out[15]~104_combout ),
	.datac(\io_out[1]~10_combout ),
	.datad(\cycleh[15]~q ),
	.cin(gnd),
	.combout(\io_out[15]~105_combout ),
	.cout());
defparam \io_out[15]~105 .lut_mask = 16'hFEEE;
defparam \io_out[15]~105 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[15]~106 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[15]~q ),
	.datad(\timeh[15]~q ),
	.cin(gnd),
	.combout(\io_out[15]~106_combout ),
	.cout());
defparam \io_out[15]~106 .lut_mask = 16'hEAC0;
defparam \io_out[15]~106 .sum_lutc_input = "datac";

dffeas \mscratch[16] (
	.clk(clock),
	.d(\_T_244[16]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[16]~q ),
	.prn(vcc));
defparam \mscratch[16] .is_wysiwyg = "true";
defparam \mscratch[16] .power_up = "low";

cyclone10lp_lcell_comb \io_out[16]~108 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[16]~q ),
	.datad(\mscratch[16]~q ),
	.cin(gnd),
	.combout(\io_out[16]~108_combout ),
	.cout());
defparam \io_out[16]~108 .lut_mask = 16'hEAC0;
defparam \io_out[16]~108 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[16]~109 (
	.dataa(ex_csr_addr_0),
	.datab(\Equal25~4_combout ),
	.datac(mepc_16),
	.datad(ex_csr_addr_1),
	.cin(gnd),
	.combout(\io_out[16]~109_combout ),
	.cout());
defparam \io_out[16]~109 .lut_mask = 16'h0080;
defparam \io_out[16]~109 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[16]~110 (
	.dataa(\io_out[16]~108_combout ),
	.datab(\io_out[16]~109_combout ),
	.datac(\io_out[1]~4_combout ),
	.datad(\time_[16]~q ),
	.cin(gnd),
	.combout(\io_out[16]~110_combout ),
	.cout());
defparam \io_out[16]~110 .lut_mask = 16'hFEEE;
defparam \io_out[16]~110 .sum_lutc_input = "datac";

dffeas \mbadaddr[16] (
	.clk(clock),
	.d(\_T_244[16]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[16]~q ),
	.prn(vcc));
defparam \mbadaddr[16] .is_wysiwyg = "true";
defparam \mbadaddr[16] .power_up = "low";

cyclone10lp_lcell_comb \io_out[16]~111 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[16]~q ),
	.datad(\mbadaddr[16]~q ),
	.cin(gnd),
	.combout(\io_out[16]~111_combout ),
	.cout());
defparam \io_out[16]~111 .lut_mask = 16'hEAC0;
defparam \io_out[16]~111 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[16]~112 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_16),
	.datad(\cycleh[16]~q ),
	.cin(gnd),
	.combout(\io_out[16]~112_combout ),
	.cout());
defparam \io_out[16]~112 .lut_mask = 16'hEAC0;
defparam \io_out[16]~112 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[16]~113 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[16]~q ),
	.datad(\timeh[16]~q ),
	.cin(gnd),
	.combout(\io_out[16]~113_combout ),
	.cout());
defparam \io_out[16]~113 .lut_mask = 16'hEAC0;
defparam \io_out[16]~113 .sum_lutc_input = "datac";

dffeas \mscratch[17] (
	.clk(clock),
	.d(\_T_244[17]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[17]~q ),
	.prn(vcc));
defparam \mscratch[17] .is_wysiwyg = "true";
defparam \mscratch[17] .power_up = "low";

cyclone10lp_lcell_comb \io_out[17]~115 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[17]~q ),
	.datad(\mscratch[17]~q ),
	.cin(gnd),
	.combout(\io_out[17]~115_combout ),
	.cout());
defparam \io_out[17]~115 .lut_mask = 16'hEAC0;
defparam \io_out[17]~115 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[17]~116 (
	.dataa(ex_csr_addr_0),
	.datab(\Equal25~4_combout ),
	.datac(mepc_17),
	.datad(ex_csr_addr_1),
	.cin(gnd),
	.combout(\io_out[17]~116_combout ),
	.cout());
defparam \io_out[17]~116 .lut_mask = 16'h0080;
defparam \io_out[17]~116 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[17]~117 (
	.dataa(\io_out[17]~115_combout ),
	.datab(\io_out[17]~116_combout ),
	.datac(\io_out[1]~4_combout ),
	.datad(\time_[17]~q ),
	.cin(gnd),
	.combout(\io_out[17]~117_combout ),
	.cout());
defparam \io_out[17]~117 .lut_mask = 16'hFEEE;
defparam \io_out[17]~117 .sum_lutc_input = "datac";

dffeas \mbadaddr[17] (
	.clk(clock),
	.d(\_T_244[17]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[17]~q ),
	.prn(vcc));
defparam \mbadaddr[17] .is_wysiwyg = "true";
defparam \mbadaddr[17] .power_up = "low";

cyclone10lp_lcell_comb \io_out[17]~118 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[17]~q ),
	.datad(\mbadaddr[17]~q ),
	.cin(gnd),
	.combout(\io_out[17]~118_combout ),
	.cout());
defparam \io_out[17]~118 .lut_mask = 16'hEAC0;
defparam \io_out[17]~118 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[17]~119 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_17),
	.datad(\cycleh[17]~q ),
	.cin(gnd),
	.combout(\io_out[17]~119_combout ),
	.cout());
defparam \io_out[17]~119 .lut_mask = 16'hEAC0;
defparam \io_out[17]~119 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[17]~120 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[17]~q ),
	.datad(\timeh[17]~q ),
	.cin(gnd),
	.combout(\io_out[17]~120_combout ),
	.cout());
defparam \io_out[17]~120 .lut_mask = 16'hEAC0;
defparam \io_out[17]~120 .sum_lutc_input = "datac";

dffeas \mscratch[18] (
	.clk(clock),
	.d(\_T_244[18]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[18]~q ),
	.prn(vcc));
defparam \mscratch[18] .is_wysiwyg = "true";
defparam \mscratch[18] .power_up = "low";

cyclone10lp_lcell_comb \io_out[18]~122 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[18]~q ),
	.datad(\mscratch[18]~q ),
	.cin(gnd),
	.combout(\io_out[18]~122_combout ),
	.cout());
defparam \io_out[18]~122 .lut_mask = 16'hEAC0;
defparam \io_out[18]~122 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[18]~123 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_18),
	.datad(\time_[18]~q ),
	.cin(gnd),
	.combout(\io_out[18]~123_combout ),
	.cout());
defparam \io_out[18]~123 .lut_mask = 16'hEAC0;
defparam \io_out[18]~123 .sum_lutc_input = "datac";

dffeas \mbadaddr[18] (
	.clk(clock),
	.d(\_T_244[18]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[18]~q ),
	.prn(vcc));
defparam \mbadaddr[18] .is_wysiwyg = "true";
defparam \mbadaddr[18] .power_up = "low";

cyclone10lp_lcell_comb \io_out[18]~124 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[18]~q ),
	.datad(\mbadaddr[18]~q ),
	.cin(gnd),
	.combout(\io_out[18]~124_combout ),
	.cout());
defparam \io_out[18]~124 .lut_mask = 16'hEAC0;
defparam \io_out[18]~124 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[18]~125 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_18),
	.datad(\cycleh[18]~q ),
	.cin(gnd),
	.combout(\io_out[18]~125_combout ),
	.cout());
defparam \io_out[18]~125 .lut_mask = 16'hEAC0;
defparam \io_out[18]~125 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[18]~126 (
	.dataa(\io_out[18]~122_combout ),
	.datab(\io_out[18]~123_combout ),
	.datac(\io_out[18]~124_combout ),
	.datad(\io_out[18]~125_combout ),
	.cin(gnd),
	.combout(\io_out[18]~126_combout ),
	.cout());
defparam \io_out[18]~126 .lut_mask = 16'hFFFE;
defparam \io_out[18]~126 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[18]~127 (
	.dataa(\io_out[1]~14_combout ),
	.datab(\instreth[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[18]~127_combout ),
	.cout());
defparam \io_out[18]~127 .lut_mask = 16'h8888;
defparam \io_out[18]~127 .sum_lutc_input = "datac";

dffeas \mscratch[19] (
	.clk(clock),
	.d(\_T_244[19]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[19]~q ),
	.prn(vcc));
defparam \mscratch[19] .is_wysiwyg = "true";
defparam \mscratch[19] .power_up = "low";

cyclone10lp_lcell_comb \io_out[19]~129 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[19]~q ),
	.datad(\mscratch[19]~q ),
	.cin(gnd),
	.combout(\io_out[19]~129_combout ),
	.cout());
defparam \io_out[19]~129 .lut_mask = 16'hEAC0;
defparam \io_out[19]~129 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[19]~130 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_19),
	.datad(\time_[19]~q ),
	.cin(gnd),
	.combout(\io_out[19]~130_combout ),
	.cout());
defparam \io_out[19]~130 .lut_mask = 16'hEAC0;
defparam \io_out[19]~130 .sum_lutc_input = "datac";

dffeas \mbadaddr[19] (
	.clk(clock),
	.d(\_T_244[19]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[19]~q ),
	.prn(vcc));
defparam \mbadaddr[19] .is_wysiwyg = "true";
defparam \mbadaddr[19] .power_up = "low";

cyclone10lp_lcell_comb \io_out[19]~131 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[19]~q ),
	.datad(\mbadaddr[19]~q ),
	.cin(gnd),
	.combout(\io_out[19]~131_combout ),
	.cout());
defparam \io_out[19]~131 .lut_mask = 16'hEAC0;
defparam \io_out[19]~131 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[19]~132 (
	.dataa(\Equal4~0_combout ),
	.datab(\Equal19~4_combout ),
	.datac(mtvec_19),
	.datad(ex_csr_addr_6),
	.cin(gnd),
	.combout(\io_out[19]~132_combout ),
	.cout());
defparam \io_out[19]~132 .lut_mask = 16'h0080;
defparam \io_out[19]~132 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[19]~133 (
	.dataa(\io_out[19]~131_combout ),
	.datab(\io_out[19]~132_combout ),
	.datac(\io_out[1]~10_combout ),
	.datad(\cycleh[19]~q ),
	.cin(gnd),
	.combout(\io_out[19]~133_combout ),
	.cout());
defparam \io_out[19]~133 .lut_mask = 16'hFEEE;
defparam \io_out[19]~133 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[19]~134 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[19]~q ),
	.datad(\timeh[19]~q ),
	.cin(gnd),
	.combout(\io_out[19]~134_combout ),
	.cout());
defparam \io_out[19]~134 .lut_mask = 16'hEAC0;
defparam \io_out[19]~134 .sum_lutc_input = "datac";

dffeas \mscratch[4] (
	.clk(clock),
	.d(\_T_244[4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[4]~q ),
	.prn(vcc));
defparam \mscratch[4] .is_wysiwyg = "true";
defparam \mscratch[4] .power_up = "low";

cyclone10lp_lcell_comb \io_out[4]~136 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[4]~q ),
	.datad(\mscratch[4]~q ),
	.cin(gnd),
	.combout(\io_out[4]~136_combout ),
	.cout());
defparam \io_out[4]~136 .lut_mask = 16'hEAC0;
defparam \io_out[4]~136 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[4]~137 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_4),
	.datad(\time_[4]~q ),
	.cin(gnd),
	.combout(\io_out[4]~137_combout ),
	.cout());
defparam \io_out[4]~137 .lut_mask = 16'hEAC0;
defparam \io_out[4]~137 .sum_lutc_input = "datac";

dffeas \mbadaddr[4] (
	.clk(clock),
	.d(\_T_244[4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[4]~q ),
	.prn(vcc));
defparam \mbadaddr[4] .is_wysiwyg = "true";
defparam \mbadaddr[4] .power_up = "low";

cyclone10lp_lcell_comb \io_out[4]~138 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[4]~q ),
	.datad(\mbadaddr[4]~q ),
	.cin(gnd),
	.combout(\io_out[4]~138_combout ),
	.cout());
defparam \io_out[4]~138 .lut_mask = 16'hEAC0;
defparam \io_out[4]~138 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \PRV1~5 (
	.dataa(io_expt1),
	.datab(isEcall),
	.datac(\_T_244[4]~1_combout ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\PRV1~5_combout ),
	.cout());
defparam \PRV1~5 .lut_mask = 16'hFDFF;
defparam \PRV1~5 .sum_lutc_input = "datac";

dffeas \PRV1[0] (
	.clk(clock),
	.d(\PRV1~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PRV1[0]~4_combout ),
	.q(\PRV1[0]~q ),
	.prn(vcc));
defparam \PRV1[0] .is_wysiwyg = "true";
defparam \PRV1[0] .power_up = "low";

cyclone10lp_lcell_comb \io_out[4]~139 (
	.dataa(\Equal19~3_combout ),
	.datab(\Equal30~0_combout ),
	.datac(\PRV1[0]~q ),
	.datad(mtvec_4),
	.cin(gnd),
	.combout(\io_out[4]~139_combout ),
	.cout());
defparam \io_out[4]~139 .lut_mask = 16'hEAC0;
defparam \io_out[4]~139 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[4]~140 (
	.dataa(\io_out[4]~138_combout ),
	.datab(\io_out[4]~139_combout ),
	.datac(\io_out[1]~10_combout ),
	.datad(\cycleh[4]~q ),
	.cin(gnd),
	.combout(\io_out[4]~140_combout ),
	.cout());
defparam \io_out[4]~140 .lut_mask = 16'hFEEE;
defparam \io_out[4]~140 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[4]~141 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[4]~q ),
	.datad(\timeh[4]~q ),
	.cin(gnd),
	.combout(\io_out[4]~141_combout ),
	.cout());
defparam \io_out[4]~141 .lut_mask = 16'hEAC0;
defparam \io_out[4]~141 .sum_lutc_input = "datac";

dffeas \mscratch[2] (
	.clk(clock),
	.d(\_T_246[2]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[2]~q ),
	.prn(vcc));
defparam \mscratch[2] .is_wysiwyg = "true";
defparam \mscratch[2] .power_up = "low";

cyclone10lp_lcell_comb \io_out[2]~143 (
	.dataa(\Equal30~0_combout ),
	.datab(\Equal25~3_combout ),
	.datac(\mscratch[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[2]~143_combout ),
	.cout());
defparam \io_out[2]~143 .lut_mask = 16'hEAEA;
defparam \io_out[2]~143 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[2]~144 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_2),
	.datad(\time_[2]~q ),
	.cin(gnd),
	.combout(\io_out[2]~144_combout ),
	.cout());
defparam \io_out[2]~144 .lut_mask = 16'hEAC0;
defparam \io_out[2]~144 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[2]~145 (
	.dataa(\io_out[2]~143_combout ),
	.datab(\io_out[2]~144_combout ),
	.datac(\io_out[1]~6_combout ),
	.datad(\cycle[2]~q ),
	.cin(gnd),
	.combout(\io_out[2]~145_combout ),
	.cout());
defparam \io_out[2]~145 .lut_mask = 16'hFEEE;
defparam \io_out[2]~145 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mcause~14 (
	.dataa(\saddrInvalid~1_combout ),
	.datab(\mcause~4_combout ),
	.datac(isEcall),
	.datad(\mcause[2]~7_combout ),
	.cin(gnd),
	.combout(\mcause~14_combout ),
	.cout());
defparam \mcause~14 .lut_mask = 16'hAA0C;
defparam \mcause~14 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mcause~15 (
	.dataa(io_expt1),
	.datab(isEcall),
	.datac(\_T_246[2]~6_combout ),
	.datad(\mcause~14_combout ),
	.cin(gnd),
	.combout(\mcause~15_combout ),
	.cout());
defparam \mcause~15 .lut_mask = 16'hFD20;
defparam \mcause~15 .sum_lutc_input = "datac";

dffeas \mcause[2] (
	.clk(clock),
	.d(\mcause~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mcause[0]~11_combout ),
	.q(\mcause[2]~q ),
	.prn(vcc));
defparam \mcause[2] .is_wysiwyg = "true";
defparam \mcause[2] .power_up = "low";

cyclone10lp_lcell_comb \io_out[2]~146 (
	.dataa(\Equal27~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[2]~q ),
	.datad(\mcause[2]~q ),
	.cin(gnd),
	.combout(\io_out[2]~146_combout ),
	.cout());
defparam \io_out[2]~146 .lut_mask = 16'hEAC0;
defparam \io_out[2]~146 .sum_lutc_input = "datac";

dffeas \mbadaddr[2] (
	.clk(clock),
	.d(\_T_246[2]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[2]~q ),
	.prn(vcc));
defparam \mbadaddr[2] .is_wysiwyg = "true";
defparam \mbadaddr[2] .power_up = "low";

cyclone10lp_lcell_comb \io_out[2]~147 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~10_combout ),
	.datac(\cycleh[2]~q ),
	.datad(\mbadaddr[2]~q ),
	.cin(gnd),
	.combout(\io_out[2]~147_combout ),
	.cout());
defparam \io_out[2]~147 .lut_mask = 16'hEAC0;
defparam \io_out[2]~147 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[2]~148 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_2),
	.datad(\timeh[2]~q ),
	.cin(gnd),
	.combout(\io_out[2]~148_combout ),
	.cout());
defparam \io_out[2]~148 .lut_mask = 16'hEAC0;
defparam \io_out[2]~148 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[2]~149 (
	.dataa(\io_out[2]~148_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[2]~149_combout ),
	.cout());
defparam \io_out[2]~149 .lut_mask = 16'hEAEA;
defparam \io_out[2]~149 .sum_lutc_input = "datac";

dffeas MSIE(
	.clk(clock),
	.d(\mtvec~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MTIE~0_combout ),
	.q(\MSIE~q ),
	.prn(vcc));
defparam MSIE.is_wysiwyg = "true";
defparam MSIE.power_up = "low";

cyclone10lp_lcell_comb \io_out[3]~151 (
	.dataa(\Equal19~3_combout ),
	.datab(\Equal21~2_combout ),
	.datac(\MSIE~q ),
	.datad(mtvec_3),
	.cin(gnd),
	.combout(\io_out[3]~151_combout ),
	.cout());
defparam \io_out[3]~151 .lut_mask = 16'hEAC0;
defparam \io_out[3]~151 .sum_lutc_input = "datac";

dffeas \mscratch[3] (
	.clk(clock),
	.d(\_T_246[3]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[3]~q ),
	.prn(vcc));
defparam \mscratch[3] .is_wysiwyg = "true";
defparam \mscratch[3] .power_up = "low";

cyclone10lp_lcell_comb \io_out[3]~152 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~12_combout ),
	.datac(\timeh[3]~q ),
	.datad(\mscratch[3]~q ),
	.cin(gnd),
	.combout(\io_out[3]~152_combout ),
	.cout());
defparam \io_out[3]~152 .lut_mask = 16'hEAC0;
defparam \io_out[3]~152 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[3]~153 (
	.dataa(\io_out[3]~151_combout ),
	.datab(\io_out[3]~152_combout ),
	.datac(\io_out[1]~4_combout ),
	.datad(\time_[3]~q ),
	.cin(gnd),
	.combout(\io_out[3]~153_combout ),
	.cout());
defparam \io_out[3]~153 .lut_mask = 16'hFEEE;
defparam \io_out[3]~153 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[3]~154 (
	.dataa(\Equal26~0_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[3]~q ),
	.datad(mepc_3),
	.cin(gnd),
	.combout(\io_out[3]~154_combout ),
	.cout());
defparam \io_out[3]~154 .lut_mask = 16'hEAC0;
defparam \io_out[3]~154 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \mcause[3]~16 (
	.dataa(io_expt1),
	.datab(isEcall),
	.datac(\_T_246[3]~8_combout ),
	.datad(ex_csr_addr_0),
	.cin(gnd),
	.combout(\mcause[3]~16_combout ),
	.cout());
defparam \mcause[3]~16 .lut_mask = 16'h20EC;
defparam \mcause[3]~16 .sum_lutc_input = "datac";

dffeas \mcause[3] (
	.clk(clock),
	.d(\mcause[3]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mcause[0]~11_combout ),
	.q(\mcause[3]~q ),
	.prn(vcc));
defparam \mcause[3] .is_wysiwyg = "true";
defparam \mcause[3] .power_up = "low";

cyclone10lp_lcell_comb \io_out[3]~155 (
	.dataa(\Equal27~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[3]~q ),
	.datad(\mcause[3]~q ),
	.cin(gnd),
	.combout(\io_out[3]~155_combout ),
	.cout());
defparam \io_out[3]~155 .lut_mask = 16'hEAC0;
defparam \io_out[3]~155 .sum_lutc_input = "datac";

dffeas \mbadaddr[3] (
	.clk(clock),
	.d(\_T_246[3]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[3]~q ),
	.prn(vcc));
defparam \mbadaddr[3] .is_wysiwyg = "true";
defparam \mbadaddr[3] .power_up = "low";

cyclone10lp_lcell_comb \io_out[3]~156 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~10_combout ),
	.datac(\cycleh[3]~q ),
	.datad(\mbadaddr[3]~q ),
	.cin(gnd),
	.combout(\io_out[3]~156_combout ),
	.cout());
defparam \io_out[3]~156 .lut_mask = 16'hEAC0;
defparam \io_out[3]~156 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MTIP~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(gnd),
	.datac(\instreth~32_combout ),
	.datad(\Equal29~2_combout ),
	.cin(gnd),
	.combout(\MTIP~0_combout ),
	.cout());
defparam \MTIP~0 .lut_mask = 16'hF555;
defparam \MTIP~0 .sum_lutc_input = "datac";

dffeas MSIP(
	.clk(clock),
	.d(\mtvec~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MTIP~0_combout ),
	.q(\MSIP~q ),
	.prn(vcc));
defparam MSIP.is_wysiwyg = "true";
defparam MSIP.power_up = "low";

cyclone10lp_lcell_comb \IE1~1 (
	.dataa(io_expt2),
	.datab(\Equal30~0_combout ),
	.datac(\wen~combout ),
	.datad(\_T_246[3]~8_combout ),
	.cin(gnd),
	.combout(\IE1~1_combout ),
	.cout());
defparam \IE1~1 .lut_mask = 16'h8000;
defparam \IE1~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \IE1~2 (
	.dataa(mcause_0),
	.datab(\IE1~1_combout ),
	.datac(\IE~q ),
	.datad(io_expt2),
	.cin(gnd),
	.combout(\IE1~2_combout ),
	.cout());
defparam \IE1~2 .lut_mask = 16'h88A8;
defparam \IE1~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \IE1~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\IE1~2_combout ),
	.datac(\IE1~0_combout ),
	.datad(\IE1~q ),
	.cin(gnd),
	.combout(\IE1~3_combout ),
	.cout());
defparam \IE1~3 .lut_mask = 16'hA888;
defparam \IE1~3 .sum_lutc_input = "datac";

dffeas IE1(
	.clk(clock),
	.d(\IE1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\IE1~q ),
	.prn(vcc));
defparam IE1.is_wysiwyg = "true";
defparam IE1.power_up = "low";

cyclone10lp_lcell_comb \io_out[3]~157 (
	.dataa(\Equal30~0_combout ),
	.datab(\Equal29~2_combout ),
	.datac(\MSIP~q ),
	.datad(\IE1~q ),
	.cin(gnd),
	.combout(\io_out[3]~157_combout ),
	.cout());
defparam \io_out[3]~157 .lut_mask = 16'hEAC0;
defparam \io_out[3]~157 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[3]~158 (
	.dataa(\io_out[3]~156_combout ),
	.datab(\io_out[3]~157_combout ),
	.datac(\io_out[1]~14_combout ),
	.datad(\instreth[3]~q ),
	.cin(gnd),
	.combout(\io_out[3]~158_combout ),
	.cout());
defparam \io_out[3]~158 .lut_mask = 16'hFEEE;
defparam \io_out[3]~158 .sum_lutc_input = "datac";

dffeas \mscratch[5] (
	.clk(clock),
	.d(\_T_244[5]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[5]~q ),
	.prn(vcc));
defparam \mscratch[5] .is_wysiwyg = "true";
defparam \mscratch[5] .power_up = "low";

cyclone10lp_lcell_comb \io_out[5]~160 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[5]~q ),
	.datad(\mscratch[5]~q ),
	.cin(gnd),
	.combout(\io_out[5]~160_combout ),
	.cout());
defparam \io_out[5]~160 .lut_mask = 16'hEAC0;
defparam \io_out[5]~160 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[5]~161 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_5),
	.datad(\time_[5]~q ),
	.cin(gnd),
	.combout(\io_out[5]~161_combout ),
	.cout());
defparam \io_out[5]~161 .lut_mask = 16'hEAC0;
defparam \io_out[5]~161 .sum_lutc_input = "datac";

dffeas \mbadaddr[5] (
	.clk(clock),
	.d(\_T_244[5]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[5]~q ),
	.prn(vcc));
defparam \mbadaddr[5] .is_wysiwyg = "true";
defparam \mbadaddr[5] .power_up = "low";

cyclone10lp_lcell_comb \io_out[5]~162 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[5]~q ),
	.datad(\mbadaddr[5]~q ),
	.cin(gnd),
	.combout(\io_out[5]~162_combout ),
	.cout());
defparam \io_out[5]~162 .lut_mask = 16'hEAC0;
defparam \io_out[5]~162 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \PRV1~6 (
	.dataa(io_expt1),
	.datab(isEcall),
	.datac(\_T_244[5]~3_combout ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\PRV1~6_combout ),
	.cout());
defparam \PRV1~6 .lut_mask = 16'hFDFF;
defparam \PRV1~6 .sum_lutc_input = "datac";

dffeas \PRV1[1] (
	.clk(clock),
	.d(\PRV1~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PRV1[0]~4_combout ),
	.q(\PRV1[1]~q ),
	.prn(vcc));
defparam \PRV1[1] .is_wysiwyg = "true";
defparam \PRV1[1] .power_up = "low";

cyclone10lp_lcell_comb \io_out[5]~163 (
	.dataa(\Equal19~3_combout ),
	.datab(\Equal30~0_combout ),
	.datac(\PRV1[1]~q ),
	.datad(mtvec_5),
	.cin(gnd),
	.combout(\io_out[5]~163_combout ),
	.cout());
defparam \io_out[5]~163 .lut_mask = 16'hEAC0;
defparam \io_out[5]~163 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[5]~164 (
	.dataa(\io_out[5]~162_combout ),
	.datab(\io_out[5]~163_combout ),
	.datac(\io_out[1]~10_combout ),
	.datad(\cycleh[5]~q ),
	.cin(gnd),
	.combout(\io_out[5]~164_combout ),
	.cout());
defparam \io_out[5]~164 .lut_mask = 16'hFEEE;
defparam \io_out[5]~164 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[5]~165 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[5]~q ),
	.datad(\timeh[5]~q ),
	.cin(gnd),
	.combout(\io_out[5]~165_combout ),
	.cout());
defparam \io_out[5]~165 .lut_mask = 16'hEAC0;
defparam \io_out[5]~165 .sum_lutc_input = "datac";

dffeas \mscratch[6] (
	.clk(clock),
	.d(\_T_244[6]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[6]~q ),
	.prn(vcc));
defparam \mscratch[6] .is_wysiwyg = "true";
defparam \mscratch[6] .power_up = "low";

cyclone10lp_lcell_comb \io_out[6]~167 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[6]~q ),
	.datad(\mscratch[6]~q ),
	.cin(gnd),
	.combout(\io_out[6]~167_combout ),
	.cout());
defparam \io_out[6]~167 .lut_mask = 16'hEAC0;
defparam \io_out[6]~167 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[6]~168 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_6),
	.datad(\time_[6]~q ),
	.cin(gnd),
	.combout(\io_out[6]~168_combout ),
	.cout());
defparam \io_out[6]~168 .lut_mask = 16'hEAC0;
defparam \io_out[6]~168 .sum_lutc_input = "datac";

dffeas \mbadaddr[6] (
	.clk(clock),
	.d(\_T_244[6]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[6]~q ),
	.prn(vcc));
defparam \mbadaddr[6] .is_wysiwyg = "true";
defparam \mbadaddr[6] .power_up = "low";

cyclone10lp_lcell_comb \io_out[6]~169 (
	.dataa(ex_csr_addr_0),
	.datab(ex_csr_addr_1),
	.datac(\Equal25~4_combout ),
	.datad(\mbadaddr[6]~q ),
	.cin(gnd),
	.combout(\io_out[6]~169_combout ),
	.cout());
defparam \io_out[6]~169 .lut_mask = 16'h8000;
defparam \io_out[6]~169 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[6]~170 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_6),
	.datad(\cycleh[6]~q ),
	.cin(gnd),
	.combout(\io_out[6]~170_combout ),
	.cout());
defparam \io_out[6]~170 .lut_mask = 16'hEAC0;
defparam \io_out[6]~170 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[6]~171 (
	.dataa(\io_out[6]~169_combout ),
	.datab(\io_out[6]~170_combout ),
	.datac(\io_out[1]~8_combout ),
	.datad(\instret[6]~q ),
	.cin(gnd),
	.combout(\io_out[6]~171_combout ),
	.cout());
defparam \io_out[6]~171 .lut_mask = 16'hFEEE;
defparam \io_out[6]~171 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[6]~172 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[6]~q ),
	.datad(\timeh[6]~q ),
	.cin(gnd),
	.combout(\io_out[6]~172_combout ),
	.cout());
defparam \io_out[6]~172 .lut_mask = 16'hEAC0;
defparam \io_out[6]~172 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \MTIE~1 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\_T_244[7]~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\MTIE~1_combout ),
	.cout());
defparam \MTIE~1 .lut_mask = 16'h8888;
defparam \MTIE~1 .sum_lutc_input = "datac";

dffeas MTIE(
	.clk(clock),
	.d(\MTIE~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MTIE~0_combout ),
	.q(\MTIE~q ),
	.prn(vcc));
defparam MTIE.is_wysiwyg = "true";
defparam MTIE.power_up = "low";

cyclone10lp_lcell_comb \io_out[7]~174 (
	.dataa(\Equal19~3_combout ),
	.datab(\Equal21~2_combout ),
	.datac(\MTIE~q ),
	.datad(mtvec_7),
	.cin(gnd),
	.combout(\io_out[7]~174_combout ),
	.cout());
defparam \io_out[7]~174 .lut_mask = 16'hEAC0;
defparam \io_out[7]~174 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[7]~175 (
	.dataa(\io_out[7]~174_combout ),
	.datab(\io_out[1]~4_combout ),
	.datac(\time_[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[7]~175_combout ),
	.cout());
defparam \io_out[7]~175 .lut_mask = 16'hEAEA;
defparam \io_out[7]~175 .sum_lutc_input = "datac";

dffeas \mscratch[7] (
	.clk(clock),
	.d(\_T_244[7]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[7]~q ),
	.prn(vcc));
defparam \mscratch[7] .is_wysiwyg = "true";
defparam \mscratch[7] .power_up = "low";

cyclone10lp_lcell_comb \io_out[7]~176 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~12_combout ),
	.datac(\timeh[7]~q ),
	.datad(\mscratch[7]~q ),
	.cin(gnd),
	.combout(\io_out[7]~176_combout ),
	.cout());
defparam \io_out[7]~176 .lut_mask = 16'hEAC0;
defparam \io_out[7]~176 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[7]~177 (
	.dataa(\Equal26~0_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[7]~q ),
	.datad(mepc_7),
	.cin(gnd),
	.combout(\io_out[7]~177_combout ),
	.cout());
defparam \io_out[7]~177 .lut_mask = 16'hEAC0;
defparam \io_out[7]~177 .sum_lutc_input = "datac";

dffeas \mbadaddr[7] (
	.clk(clock),
	.d(\_T_244[7]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[7]~q ),
	.prn(vcc));
defparam \mbadaddr[7] .is_wysiwyg = "true";
defparam \mbadaddr[7] .power_up = "low";

cyclone10lp_lcell_comb \io_out[7]~178 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[7]~q ),
	.datad(\mbadaddr[7]~q ),
	.cin(gnd),
	.combout(\io_out[7]~178_combout ),
	.cout());
defparam \io_out[7]~178 .lut_mask = 16'hEAC0;
defparam \io_out[7]~178 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[7]~179 (
	.dataa(\io_out[7]~175_combout ),
	.datab(\io_out[7]~176_combout ),
	.datac(\io_out[7]~177_combout ),
	.datad(\io_out[7]~178_combout ),
	.cin(gnd),
	.combout(\io_out[7]~179_combout ),
	.cout());
defparam \io_out[7]~179 .lut_mask = 16'hFFFE;
defparam \io_out[7]~179 .sum_lutc_input = "datac";

dffeas MTIP(
	.clk(clock),
	.d(\MTIE~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MTIP~0_combout ),
	.q(\MTIP~q ),
	.prn(vcc));
defparam MTIP.is_wysiwyg = "true";
defparam MTIP.power_up = "low";

cyclone10lp_lcell_comb \io_out[7]~180 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal29~2_combout ),
	.datac(\MTIP~q ),
	.datad(\cycleh[7]~q ),
	.cin(gnd),
	.combout(\io_out[7]~180_combout ),
	.cout());
defparam \io_out[7]~180 .lut_mask = 16'hEAC0;
defparam \io_out[7]~180 .sum_lutc_input = "datac";

dffeas \mscratch[20] (
	.clk(clock),
	.d(\_T_244[20]~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[20]~q ),
	.prn(vcc));
defparam \mscratch[20] .is_wysiwyg = "true";
defparam \mscratch[20] .power_up = "low";

cyclone10lp_lcell_comb \io_out[20]~182 (
	.dataa(\Equal16~2_combout ),
	.datab(\Equal25~3_combout ),
	.datac(\mscratch[20]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[20]~182_combout ),
	.cout());
defparam \io_out[20]~182 .lut_mask = 16'hEAEA;
defparam \io_out[20]~182 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[20]~183 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_20),
	.datad(\time_[20]~q ),
	.cin(gnd),
	.combout(\io_out[20]~183_combout ),
	.cout());
defparam \io_out[20]~183 .lut_mask = 16'hEAC0;
defparam \io_out[20]~183 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[20]~184 (
	.dataa(\io_out[20]~182_combout ),
	.datab(\io_out[20]~183_combout ),
	.datac(\io_out[1]~6_combout ),
	.datad(\cycle[20]~q ),
	.cin(gnd),
	.combout(\io_out[20]~184_combout ),
	.cout());
defparam \io_out[20]~184 .lut_mask = 16'hFEEE;
defparam \io_out[20]~184 .sum_lutc_input = "datac";

dffeas \mbadaddr[20] (
	.clk(clock),
	.d(\_T_244[20]~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[20]~q ),
	.prn(vcc));
defparam \mbadaddr[20] .is_wysiwyg = "true";
defparam \mbadaddr[20] .power_up = "low";

cyclone10lp_lcell_comb \io_out[20]~185 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[20]~q ),
	.datad(\mbadaddr[20]~q ),
	.cin(gnd),
	.combout(\io_out[20]~185_combout ),
	.cout());
defparam \io_out[20]~185 .lut_mask = 16'hEAC0;
defparam \io_out[20]~185 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[20]~186 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_20),
	.datad(\cycleh[20]~q ),
	.cin(gnd),
	.combout(\io_out[20]~186_combout ),
	.cout());
defparam \io_out[20]~186 .lut_mask = 16'hEAC0;
defparam \io_out[20]~186 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[20]~187 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[20]~q ),
	.datad(\timeh[20]~q ),
	.cin(gnd),
	.combout(\io_out[20]~187_combout ),
	.cout());
defparam \io_out[20]~187 .lut_mask = 16'hEAC0;
defparam \io_out[20]~187 .sum_lutc_input = "datac";

dffeas \mscratch[21] (
	.clk(clock),
	.d(\_T_244[21]~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[21]~q ),
	.prn(vcc));
defparam \mscratch[21] .is_wysiwyg = "true";
defparam \mscratch[21] .power_up = "low";

cyclone10lp_lcell_comb \io_out[21]~189 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[21]~q ),
	.datad(\mscratch[21]~q ),
	.cin(gnd),
	.combout(\io_out[21]~189_combout ),
	.cout());
defparam \io_out[21]~189 .lut_mask = 16'hEAC0;
defparam \io_out[21]~189 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[21]~190 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_21),
	.datad(\time_[21]~q ),
	.cin(gnd),
	.combout(\io_out[21]~190_combout ),
	.cout());
defparam \io_out[21]~190 .lut_mask = 16'hEAC0;
defparam \io_out[21]~190 .sum_lutc_input = "datac";

dffeas \mbadaddr[21] (
	.clk(clock),
	.d(\_T_244[21]~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[21]~q ),
	.prn(vcc));
defparam \mbadaddr[21] .is_wysiwyg = "true";
defparam \mbadaddr[21] .power_up = "low";

cyclone10lp_lcell_comb \io_out[21]~191 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[21]~q ),
	.datad(\mbadaddr[21]~q ),
	.cin(gnd),
	.combout(\io_out[21]~191_combout ),
	.cout());
defparam \io_out[21]~191 .lut_mask = 16'hEAC0;
defparam \io_out[21]~191 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[21]~192 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_21),
	.datad(\cycleh[21]~q ),
	.cin(gnd),
	.combout(\io_out[21]~192_combout ),
	.cout());
defparam \io_out[21]~192 .lut_mask = 16'hEAC0;
defparam \io_out[21]~192 .sum_lutc_input = "datac";

dffeas \mscratch[22] (
	.clk(clock),
	.d(\_T_244[22]~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[22]~q ),
	.prn(vcc));
defparam \mscratch[22] .is_wysiwyg = "true";
defparam \mscratch[22] .power_up = "low";

cyclone10lp_lcell_comb \io_out[22]~196 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[22]~q ),
	.datad(\mscratch[22]~q ),
	.cin(gnd),
	.combout(\io_out[22]~196_combout ),
	.cout());
defparam \io_out[22]~196 .lut_mask = 16'hEAC0;
defparam \io_out[22]~196 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[22]~197 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_22),
	.datad(\time_[22]~q ),
	.cin(gnd),
	.combout(\io_out[22]~197_combout ),
	.cout());
defparam \io_out[22]~197 .lut_mask = 16'hEAC0;
defparam \io_out[22]~197 .sum_lutc_input = "datac";

dffeas \mbadaddr[22] (
	.clk(clock),
	.d(\_T_244[22]~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[22]~q ),
	.prn(vcc));
defparam \mbadaddr[22] .is_wysiwyg = "true";
defparam \mbadaddr[22] .power_up = "low";

cyclone10lp_lcell_comb \io_out[22]~198 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[22]~q ),
	.datad(\mbadaddr[22]~q ),
	.cin(gnd),
	.combout(\io_out[22]~198_combout ),
	.cout());
defparam \io_out[22]~198 .lut_mask = 16'hEAC0;
defparam \io_out[22]~198 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[22]~199 (
	.dataa(\Equal19~2_combout ),
	.datab(\Equal19~4_combout ),
	.datac(mtvec_22),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[22]~199_combout ),
	.cout());
defparam \io_out[22]~199 .lut_mask = 16'h8080;
defparam \io_out[22]~199 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[22]~200 (
	.dataa(\io_out[22]~198_combout ),
	.datab(\io_out[22]~199_combout ),
	.datac(\io_out[1]~10_combout ),
	.datad(\cycleh[22]~q ),
	.cin(gnd),
	.combout(\io_out[22]~200_combout ),
	.cout());
defparam \io_out[22]~200 .lut_mask = 16'hFEEE;
defparam \io_out[22]~200 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[22]~201 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[22]~q ),
	.datad(\timeh[22]~q ),
	.cin(gnd),
	.combout(\io_out[22]~201_combout ),
	.cout());
defparam \io_out[22]~201 .lut_mask = 16'hEAC0;
defparam \io_out[22]~201 .sum_lutc_input = "datac";

dffeas \mscratch[23] (
	.clk(clock),
	.d(\_T_244[23]~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[23]~q ),
	.prn(vcc));
defparam \mscratch[23] .is_wysiwyg = "true";
defparam \mscratch[23] .power_up = "low";

cyclone10lp_lcell_comb \io_out[23]~203 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[23]~q ),
	.datad(\mscratch[23]~q ),
	.cin(gnd),
	.combout(\io_out[23]~203_combout ),
	.cout());
defparam \io_out[23]~203 .lut_mask = 16'hEAC0;
defparam \io_out[23]~203 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[23]~204 (
	.dataa(ex_csr_addr_0),
	.datab(\Equal25~4_combout ),
	.datac(mepc_23),
	.datad(ex_csr_addr_1),
	.cin(gnd),
	.combout(\io_out[23]~204_combout ),
	.cout());
defparam \io_out[23]~204 .lut_mask = 16'h0080;
defparam \io_out[23]~204 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[23]~205 (
	.dataa(\io_out[23]~203_combout ),
	.datab(\io_out[23]~204_combout ),
	.datac(\io_out[1]~4_combout ),
	.datad(\time_[23]~q ),
	.cin(gnd),
	.combout(\io_out[23]~205_combout ),
	.cout());
defparam \io_out[23]~205 .lut_mask = 16'hFEEE;
defparam \io_out[23]~205 .sum_lutc_input = "datac";

dffeas \mbadaddr[23] (
	.clk(clock),
	.d(\_T_244[23]~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[23]~q ),
	.prn(vcc));
defparam \mbadaddr[23] .is_wysiwyg = "true";
defparam \mbadaddr[23] .power_up = "low";

cyclone10lp_lcell_comb \io_out[23]~206 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[23]~q ),
	.datad(\mbadaddr[23]~q ),
	.cin(gnd),
	.combout(\io_out[23]~206_combout ),
	.cout());
defparam \io_out[23]~206 .lut_mask = 16'hEAC0;
defparam \io_out[23]~206 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[23]~207 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_23),
	.datad(\cycleh[23]~q ),
	.cin(gnd),
	.combout(\io_out[23]~207_combout ),
	.cout());
defparam \io_out[23]~207 .lut_mask = 16'hEAC0;
defparam \io_out[23]~207 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[23]~208 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[23]~q ),
	.datad(\timeh[23]~q ),
	.cin(gnd),
	.combout(\io_out[23]~208_combout ),
	.cout());
defparam \io_out[23]~208 .lut_mask = 16'hEAC0;
defparam \io_out[23]~208 .sum_lutc_input = "datac";

dffeas \mscratch[24] (
	.clk(clock),
	.d(\_T_244[24]~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[24]~q ),
	.prn(vcc));
defparam \mscratch[24] .is_wysiwyg = "true";
defparam \mscratch[24] .power_up = "low";

cyclone10lp_lcell_comb \io_out[24]~210 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[24]~q ),
	.datad(\mscratch[24]~q ),
	.cin(gnd),
	.combout(\io_out[24]~210_combout ),
	.cout());
defparam \io_out[24]~210 .lut_mask = 16'hEAC0;
defparam \io_out[24]~210 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[24]~211 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_24),
	.datad(\time_[24]~q ),
	.cin(gnd),
	.combout(\io_out[24]~211_combout ),
	.cout());
defparam \io_out[24]~211 .lut_mask = 16'hEAC0;
defparam \io_out[24]~211 .sum_lutc_input = "datac";

dffeas \mbadaddr[24] (
	.clk(clock),
	.d(\_T_244[24]~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[24]~q ),
	.prn(vcc));
defparam \mbadaddr[24] .is_wysiwyg = "true";
defparam \mbadaddr[24] .power_up = "low";

cyclone10lp_lcell_comb \io_out[24]~212 (
	.dataa(ex_csr_addr_0),
	.datab(ex_csr_addr_1),
	.datac(\Equal25~4_combout ),
	.datad(\mbadaddr[24]~q ),
	.cin(gnd),
	.combout(\io_out[24]~212_combout ),
	.cout());
defparam \io_out[24]~212 .lut_mask = 16'h8000;
defparam \io_out[24]~212 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[24]~213 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_24),
	.datad(\cycleh[24]~q ),
	.cin(gnd),
	.combout(\io_out[24]~213_combout ),
	.cout());
defparam \io_out[24]~213 .lut_mask = 16'hEAC0;
defparam \io_out[24]~213 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[24]~214 (
	.dataa(\io_out[24]~212_combout ),
	.datab(\io_out[24]~213_combout ),
	.datac(\io_out[1]~8_combout ),
	.datad(\instret[24]~q ),
	.cin(gnd),
	.combout(\io_out[24]~214_combout ),
	.cout());
defparam \io_out[24]~214 .lut_mask = 16'hFEEE;
defparam \io_out[24]~214 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[24]~215 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[24]~q ),
	.datad(\timeh[24]~q ),
	.cin(gnd),
	.combout(\io_out[24]~215_combout ),
	.cout());
defparam \io_out[24]~215 .lut_mask = 16'hEAC0;
defparam \io_out[24]~215 .sum_lutc_input = "datac";

dffeas \mscratch[25] (
	.clk(clock),
	.d(\_T_244[25]~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[25]~q ),
	.prn(vcc));
defparam \mscratch[25] .is_wysiwyg = "true";
defparam \mscratch[25] .power_up = "low";

cyclone10lp_lcell_comb \io_out[25]~217 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[25]~q ),
	.datad(\mscratch[25]~q ),
	.cin(gnd),
	.combout(\io_out[25]~217_combout ),
	.cout());
defparam \io_out[25]~217 .lut_mask = 16'hEAC0;
defparam \io_out[25]~217 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[25]~218 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_25),
	.datad(\time_[25]~q ),
	.cin(gnd),
	.combout(\io_out[25]~218_combout ),
	.cout());
defparam \io_out[25]~218 .lut_mask = 16'hEAC0;
defparam \io_out[25]~218 .sum_lutc_input = "datac";

dffeas \mbadaddr[25] (
	.clk(clock),
	.d(\_T_244[25]~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[25]~q ),
	.prn(vcc));
defparam \mbadaddr[25] .is_wysiwyg = "true";
defparam \mbadaddr[25] .power_up = "low";

cyclone10lp_lcell_comb \io_out[25]~219 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[25]~q ),
	.datad(\mbadaddr[25]~q ),
	.cin(gnd),
	.combout(\io_out[25]~219_combout ),
	.cout());
defparam \io_out[25]~219 .lut_mask = 16'hEAC0;
defparam \io_out[25]~219 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[25]~220 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_25),
	.datad(\cycleh[25]~q ),
	.cin(gnd),
	.combout(\io_out[25]~220_combout ),
	.cout());
defparam \io_out[25]~220 .lut_mask = 16'hEAC0;
defparam \io_out[25]~220 .sum_lutc_input = "datac";

dffeas \mscratch[26] (
	.clk(clock),
	.d(\_T_244[26]~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[26]~q ),
	.prn(vcc));
defparam \mscratch[26] .is_wysiwyg = "true";
defparam \mscratch[26] .power_up = "low";

cyclone10lp_lcell_comb \io_out[26]~224 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[26]~q ),
	.datad(\mscratch[26]~q ),
	.cin(gnd),
	.combout(\io_out[26]~224_combout ),
	.cout());
defparam \io_out[26]~224 .lut_mask = 16'hEAC0;
defparam \io_out[26]~224 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[26]~225 (
	.dataa(\Equal26~0_combout ),
	.datab(mepc_26),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\io_out[26]~225_combout ),
	.cout());
defparam \io_out[26]~225 .lut_mask = 16'h8888;
defparam \io_out[26]~225 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[26]~226 (
	.dataa(\io_out[26]~224_combout ),
	.datab(\io_out[26]~225_combout ),
	.datac(\io_out[1]~4_combout ),
	.datad(\time_[26]~q ),
	.cin(gnd),
	.combout(\io_out[26]~226_combout ),
	.cout());
defparam \io_out[26]~226 .lut_mask = 16'hFEEE;
defparam \io_out[26]~226 .sum_lutc_input = "datac";

dffeas \mbadaddr[26] (
	.clk(clock),
	.d(\_T_244[26]~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[26]~q ),
	.prn(vcc));
defparam \mbadaddr[26] .is_wysiwyg = "true";
defparam \mbadaddr[26] .power_up = "low";

cyclone10lp_lcell_comb \io_out[26]~227 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[26]~q ),
	.datad(\mbadaddr[26]~q ),
	.cin(gnd),
	.combout(\io_out[26]~227_combout ),
	.cout());
defparam \io_out[26]~227 .lut_mask = 16'hEAC0;
defparam \io_out[26]~227 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[26]~228 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_26),
	.datad(\cycleh[26]~q ),
	.cin(gnd),
	.combout(\io_out[26]~228_combout ),
	.cout());
defparam \io_out[26]~228 .lut_mask = 16'hEAC0;
defparam \io_out[26]~228 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[26]~229 (
	.dataa(\io_out[1]~12_combout ),
	.datab(\io_out[1]~14_combout ),
	.datac(\instreth[26]~q ),
	.datad(\timeh[26]~q ),
	.cin(gnd),
	.combout(\io_out[26]~229_combout ),
	.cout());
defparam \io_out[26]~229 .lut_mask = 16'hEAC0;
defparam \io_out[26]~229 .sum_lutc_input = "datac";

dffeas \mscratch[27] (
	.clk(clock),
	.d(\_T_244[27]~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mscratch[0]~0_combout ),
	.q(\mscratch[27]~q ),
	.prn(vcc));
defparam \mscratch[27] .is_wysiwyg = "true";
defparam \mscratch[27] .power_up = "low";

cyclone10lp_lcell_comb \io_out[27]~231 (
	.dataa(\Equal25~3_combout ),
	.datab(\io_out[1]~6_combout ),
	.datac(\cycle[27]~q ),
	.datad(\mscratch[27]~q ),
	.cin(gnd),
	.combout(\io_out[27]~231_combout ),
	.cout());
defparam \io_out[27]~231 .lut_mask = 16'hEAC0;
defparam \io_out[27]~231 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[27]~232 (
	.dataa(\io_out[1]~4_combout ),
	.datab(\Equal26~0_combout ),
	.datac(mepc_27),
	.datad(\time_[27]~q ),
	.cin(gnd),
	.combout(\io_out[27]~232_combout ),
	.cout());
defparam \io_out[27]~232 .lut_mask = 16'hEAC0;
defparam \io_out[27]~232 .sum_lutc_input = "datac";

dffeas \mbadaddr[27] (
	.clk(clock),
	.d(\_T_244[27]~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mbadaddr[0]~0_combout ),
	.q(\mbadaddr[27]~q ),
	.prn(vcc));
defparam \mbadaddr[27] .is_wysiwyg = "true";
defparam \mbadaddr[27] .power_up = "low";

cyclone10lp_lcell_comb \io_out[27]~233 (
	.dataa(\Equal28~0_combout ),
	.datab(\io_out[1]~8_combout ),
	.datac(\instret[27]~q ),
	.datad(\mbadaddr[27]~q ),
	.cin(gnd),
	.combout(\io_out[27]~233_combout ),
	.cout());
defparam \io_out[27]~233 .lut_mask = 16'hEAC0;
defparam \io_out[27]~233 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \io_out[27]~234 (
	.dataa(\io_out[1]~10_combout ),
	.datab(\Equal19~3_combout ),
	.datac(mtvec_27),
	.datad(\cycleh[27]~q ),
	.cin(gnd),
	.combout(\io_out[27]~234_combout ),
	.cout());
defparam \io_out[27]~234 .lut_mask = 16'hEAC0;
defparam \io_out[27]~234 .sum_lutc_input = "datac";

endmodule

module kyogenrv_fpga_kyogenrv_fpga_mm_interconnect_0 (
	av_readdata_pre_1,
	av_readdata_pre_0,
	waitrequest_reset_override,
	wait_latency_counter_0,
	mem_ctrl_mem_wr10,
	wait_latency_counter_1,
	altera_reset_synchronizer_int_chain_out,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_30,
	av_readdata_pre_31,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata_pre_18,
	av_readdata_pre_19,
	av_readdata_pre_4,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_20,
	av_readdata_pre_21,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_27,
	readdata_1,
	readdata_0,
	mem_ctrl_mem_wr00,
	mem_ctrl_mem_wr01,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	readdata_8,
	readdata_9,
	readdata_10,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_17,
	readdata_18,
	readdata_19,
	readdata_4,
	readdata_2,
	readdata_3,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_20,
	readdata_21,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_27,
	read_latency_shift_reg_0,
	clk_clk)/* synthesis synthesis_greybox=0 */;
output 	av_readdata_pre_1;
output 	av_readdata_pre_0;
output 	waitrequest_reset_override;
output 	wait_latency_counter_0;
input 	mem_ctrl_mem_wr10;
output 	wait_latency_counter_1;
input 	altera_reset_synchronizer_int_chain_out;
output 	av_readdata_pre_28;
output 	av_readdata_pre_29;
output 	av_readdata_pre_30;
output 	av_readdata_pre_31;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_16;
output 	av_readdata_pre_17;
output 	av_readdata_pre_18;
output 	av_readdata_pre_19;
output 	av_readdata_pre_4;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_20;
output 	av_readdata_pre_21;
output 	av_readdata_pre_22;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_26;
output 	av_readdata_pre_27;
input 	readdata_1;
input 	readdata_0;
input 	mem_ctrl_mem_wr00;
input 	mem_ctrl_mem_wr01;
input 	readdata_28;
input 	readdata_29;
input 	readdata_30;
input 	readdata_31;
input 	readdata_8;
input 	readdata_9;
input 	readdata_10;
input 	readdata_11;
input 	readdata_12;
input 	readdata_13;
input 	readdata_14;
input 	readdata_15;
input 	readdata_16;
input 	readdata_17;
input 	readdata_18;
input 	readdata_19;
input 	readdata_4;
input 	readdata_2;
input 	readdata_3;
input 	readdata_5;
input 	readdata_6;
input 	readdata_7;
input 	readdata_20;
input 	readdata_21;
input 	readdata_22;
input 	readdata_23;
input 	readdata_24;
input 	readdata_25;
input 	readdata_26;
input 	readdata_27;
output 	read_latency_shift_reg_0;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



kyogenrv_fpga_altera_merlin_slave_translator pio_0_s1_translator(
	.av_readdata_pre_1(av_readdata_pre_1),
	.av_readdata_pre_0(av_readdata_pre_0),
	.waitrequest_reset_override1(waitrequest_reset_override),
	.wait_latency_counter_0(wait_latency_counter_0),
	.mem_ctrl_mem_wr10(mem_ctrl_mem_wr10),
	.wait_latency_counter_1(wait_latency_counter_1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.av_readdata_pre_28(av_readdata_pre_28),
	.av_readdata_pre_29(av_readdata_pre_29),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata_pre_31(av_readdata_pre_31),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_16(av_readdata_pre_16),
	.av_readdata_pre_17(av_readdata_pre_17),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_19(av_readdata_pre_19),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_2(av_readdata_pre_2),
	.av_readdata_pre_3(av_readdata_pre_3),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_6(av_readdata_pre_6),
	.av_readdata_pre_7(av_readdata_pre_7),
	.av_readdata_pre_20(av_readdata_pre_20),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_22(av_readdata_pre_22),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_24(av_readdata_pre_24),
	.av_readdata_pre_25(av_readdata_pre_25),
	.av_readdata_pre_26(av_readdata_pre_26),
	.av_readdata_pre_27(av_readdata_pre_27),
	.av_readdata({readdata_31,readdata_30,readdata_29,readdata_28,readdata_27,readdata_26,readdata_25,readdata_24,readdata_23,readdata_22,readdata_21,readdata_20,readdata_19,readdata_18,readdata_17,readdata_16,readdata_15,readdata_14,readdata_13,readdata_12,readdata_11,readdata_10,readdata_9,
readdata_8,readdata_7,readdata_6,readdata_5,readdata_4,readdata_3,readdata_2,readdata_1,readdata_0}),
	.mem_ctrl_mem_wr00(mem_ctrl_mem_wr00),
	.mem_ctrl_mem_wr01(mem_ctrl_mem_wr01),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.clk(clk_clk));

endmodule

module kyogenrv_fpga_altera_merlin_slave_translator (
	av_readdata_pre_1,
	av_readdata_pre_0,
	waitrequest_reset_override1,
	wait_latency_counter_0,
	mem_ctrl_mem_wr10,
	wait_latency_counter_1,
	reset,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_30,
	av_readdata_pre_31,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata_pre_18,
	av_readdata_pre_19,
	av_readdata_pre_4,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_20,
	av_readdata_pre_21,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_27,
	av_readdata,
	mem_ctrl_mem_wr00,
	mem_ctrl_mem_wr01,
	read_latency_shift_reg_0,
	clk)/* synthesis synthesis_greybox=0 */;
output 	av_readdata_pre_1;
output 	av_readdata_pre_0;
output 	waitrequest_reset_override1;
output 	wait_latency_counter_0;
input 	mem_ctrl_mem_wr10;
output 	wait_latency_counter_1;
input 	reset;
output 	av_readdata_pre_28;
output 	av_readdata_pre_29;
output 	av_readdata_pre_30;
output 	av_readdata_pre_31;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_16;
output 	av_readdata_pre_17;
output 	av_readdata_pre_18;
output 	av_readdata_pre_19;
output 	av_readdata_pre_4;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_20;
output 	av_readdata_pre_21;
output 	av_readdata_pre_22;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_26;
output 	av_readdata_pre_27;
input 	[31:0] av_readdata;
input 	mem_ctrl_mem_wr00;
input 	mem_ctrl_mem_wr01;
output 	read_latency_shift_reg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~0_combout ;


dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas waitrequest_reset_override(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest_reset_override1),
	.prn(vcc));
defparam waitrequest_reset_override.is_wysiwyg = "true";
defparam waitrequest_reset_override.power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclone10lp_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(waitrequest_reset_override1),
	.datab(wait_latency_counter_1),
	.datac(wait_latency_counter_0),
	.datad(mem_ctrl_mem_wr10),
	.cin(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.cout());
defparam \wait_latency_counter[0]~0 .lut_mask = 16'hA88A;
defparam \wait_latency_counter[0]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter~1 (
	.dataa(wait_latency_counter_0),
	.datab(gnd),
	.datac(mem_ctrl_mem_wr00),
	.datad(\wait_latency_counter[0]~0_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.cout());
defparam \wait_latency_counter~1 .lut_mask = 16'h5000;
defparam \wait_latency_counter~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \wait_latency_counter~2 (
	.dataa(mem_ctrl_mem_wr00),
	.datab(\wait_latency_counter[0]~0_combout ),
	.datac(wait_latency_counter_0),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'h0880;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \read_latency_shift_reg~0 (
	.dataa(wait_latency_counter_0),
	.datab(waitrequest_reset_override1),
	.datac(mem_ctrl_mem_wr01),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'h0080;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module kyogenrv_fpga_kyogenrv_fpga_mm_interconnect_1 (
	waitrequest_reset_override,
	read_latency_shift_reg_0,
	altera_reset_synchronizer_int_chain_out,
	w_req,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
output 	read_latency_shift_reg_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	w_req;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



kyogenrv_fpga_altera_merlin_slave_translator_1 onchip_memory2_0_s1_translator(
	.waitrequest_reset_override(waitrequest_reset_override),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.reset(altera_reset_synchronizer_int_chain_out),
	.w_req(w_req),
	.clk(clk_clk));

endmodule

module kyogenrv_fpga_altera_merlin_slave_translator_1 (
	waitrequest_reset_override,
	read_latency_shift_reg_0,
	reset,
	w_req,
	clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
output 	read_latency_shift_reg_0;
input 	reset;
input 	w_req;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclone10lp_lcell_comb \read_latency_shift_reg~0 (
	.dataa(w_req),
	.datab(gnd),
	.datac(gnd),
	.datad(waitrequest_reset_override),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'h5500;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module kyogenrv_fpga_kyogenrv_fpga_onchip_memory2_0 (
	q_a_16,
	q_a_15,
	q_a_18,
	q_a_17,
	q_a_19,
	q_a_21,
	q_a_20,
	q_a_23,
	q_a_22,
	q_a_24,
	q_a_14,
	q_a_13,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	q_a_12,
	q_a_10,
	q_a_11,
	q_a_25,
	q_a_30,
	q_a_0,
	q_a_1,
	q_a_3,
	q_a_2,
	q_a_4,
	q_a_26,
	q_a_27,
	q_a_31,
	q_a_28,
	q_a_29,
	w_req,
	io_imem_add_addr_2,
	io_imem_add_addr_3,
	io_imem_add_addr_4,
	io_imem_add_addr_5,
	io_imem_add_addr_6,
	io_imem_add_addr_7,
	io_imem_add_addr_8,
	io_imem_add_addr_9,
	io_imem_add_addr_10,
	io_imem_add_addr_11,
	io_imem_add_addr_12,
	io_imem_add_addr_13,
	io_imem_add_addr_14,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=0 */;
output 	q_a_16;
output 	q_a_15;
output 	q_a_18;
output 	q_a_17;
output 	q_a_19;
output 	q_a_21;
output 	q_a_20;
output 	q_a_23;
output 	q_a_22;
output 	q_a_24;
output 	q_a_14;
output 	q_a_13;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
output 	q_a_12;
output 	q_a_10;
output 	q_a_11;
output 	q_a_25;
output 	q_a_30;
output 	q_a_0;
output 	q_a_1;
output 	q_a_3;
output 	q_a_2;
output 	q_a_4;
output 	q_a_26;
output 	q_a_27;
output 	q_a_31;
output 	q_a_28;
output 	q_a_29;
input 	w_req;
input 	io_imem_add_addr_2;
input 	io_imem_add_addr_3;
input 	io_imem_add_addr_4;
input 	io_imem_add_addr_5;
input 	io_imem_add_addr_6;
input 	io_imem_add_addr_7;
input 	io_imem_add_addr_8;
input 	io_imem_add_addr_9;
input 	io_imem_add_addr_10;
input 	io_imem_add_addr_11;
input 	io_imem_add_addr_12;
input 	io_imem_add_addr_13;
input 	io_imem_add_addr_14;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



kyogenrv_fpga_altsyncram_1 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.wren_a(w_req),
	.address_a({io_imem_add_addr_14,io_imem_add_addr_13,io_imem_add_addr_12,io_imem_add_addr_11,io_imem_add_addr_10,io_imem_add_addr_9,io_imem_add_addr_8,io_imem_add_addr_7,io_imem_add_addr_6,io_imem_add_addr_5,io_imem_add_addr_4,io_imem_add_addr_3,io_imem_add_addr_2}),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,GND_port,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.clock0(clk_clk));

endmodule

module kyogenrv_fpga_altsyncram_1 (
	q_a,
	wren_a,
	address_a,
	data_a,
	clock0)/* synthesis synthesis_greybox=0 */;
output 	[31:0] q_a;
input 	wren_a;
input 	[12:0] address_a;
input 	[31:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



kyogenrv_fpga_altsyncram_63i1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.wren_a(wren_a),
	.address_a({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.data_a({data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16],data_a[16]}),
	.clock0(clock0));

endmodule

module kyogenrv_fpga_altsyncram_63i1 (
	q_a,
	wren_a,
	address_a,
	data_a,
	clock0)/* synthesis synthesis_greybox=0 */;
output 	[31:0] q_a;
input 	wren_a;
input 	[12:0] address_a;
input 	[31:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

cyclone10lp_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 13;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 8191;
defparam ram_block1a16.port_a_logical_ram_depth = 8192;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a16.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a16.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a16.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 13;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 8191;
defparam ram_block1a15.port_a_logical_ram_depth = 8192;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a15.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a15.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a15.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000068;

cyclone10lp_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 13;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 8191;
defparam ram_block1a18.port_a_logical_ram_depth = 8192;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a18.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a18.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a18.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 13;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 8191;
defparam ram_block1a17.port_a_logical_ram_depth = 8192;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a17.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a17.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a17.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 13;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 8191;
defparam ram_block1a19.port_a_logical_ram_depth = 8192;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a19.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a19.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a19.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 13;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 8191;
defparam ram_block1a21.port_a_logical_ram_depth = 8192;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a21.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a21.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a21.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000070;

cyclone10lp_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 13;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 8191;
defparam ram_block1a20.port_a_logical_ram_depth = 8192;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a20.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a20.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a20.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 13;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 8191;
defparam ram_block1a23.port_a_logical_ram_depth = 8192;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a23.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a23.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a23.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;

cyclone10lp_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 13;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 8191;
defparam ram_block1a22.port_a_logical_ram_depth = 8192;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a22.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a22.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a22.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 13;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 8191;
defparam ram_block1a24.port_a_logical_ram_depth = 8192;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a24.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a24.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a24.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 13;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 8191;
defparam ram_block1a14.port_a_logical_ram_depth = 8192;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a14.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a14.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a14.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 13;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 8191;
defparam ram_block1a13.port_a_logical_ram_depth = 8192;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a13.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a13.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a13.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020;

cyclone10lp_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 13;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 8191;
defparam ram_block1a5.port_a_logical_ram_depth = 8192;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a5.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a5.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a5.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000E8;

cyclone10lp_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 13;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 8191;
defparam ram_block1a6.port_a_logical_ram_depth = 8192;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a6.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a6.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a6.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000080;

cyclone10lp_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 13;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 8191;
defparam ram_block1a7.port_a_logical_ram_depth = 8192;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a7.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a7.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a7.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008;

cyclone10lp_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 13;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 8191;
defparam ram_block1a8.port_a_logical_ram_depth = 8192;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a8.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a8.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a8.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;

cyclone10lp_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 13;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 8191;
defparam ram_block1a9.port_a_logical_ram_depth = 8192;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a9.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a9.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a9.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 13;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 8191;
defparam ram_block1a12.port_a_logical_ram_depth = 8192;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a12.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a12.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a12.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 13;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 8191;
defparam ram_block1a10.port_a_logical_ram_depth = 8192;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a10.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a10.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a10.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 13;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 8191;
defparam ram_block1a11.port_a_logical_ram_depth = 8192;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a11.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a11.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a11.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 13;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 8191;
defparam ram_block1a25.port_a_logical_ram_depth = 8192;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a25.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a25.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a25.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;

cyclone10lp_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 13;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 8191;
defparam ram_block1a30.port_a_logical_ram_depth = 8192;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a30.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a30.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a30.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 13;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 8191;
defparam ram_block1a0.port_a_logical_ram_depth = 8192;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a0.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a0.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a0.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF;

cyclone10lp_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 13;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 8191;
defparam ram_block1a1.port_a_logical_ram_depth = 8192;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a1.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a1.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a1.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF;

cyclone10lp_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 13;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 8191;
defparam ram_block1a3.port_a_logical_ram_depth = 8192;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a3.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a3.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a3.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000080;

cyclone10lp_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 13;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 8191;
defparam ram_block1a2.port_a_logical_ram_depth = 8192;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a2.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a2.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a2.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000088;

cyclone10lp_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 13;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 8191;
defparam ram_block1a4.port_a_logical_ram_depth = 8192;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a4.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a4.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a4.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001F;

cyclone10lp_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 13;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 8191;
defparam ram_block1a26.port_a_logical_ram_depth = 8192;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a26.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a26.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a26.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 13;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 8191;
defparam ram_block1a27.port_a_logical_ram_depth = 8192;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a27.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a27.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a27.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;

cyclone10lp_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 13;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 8191;
defparam ram_block1a31.port_a_logical_ram_depth = 8192;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a31.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a31.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a31.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 13;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 8191;
defparam ram_block1a28.port_a_logical_ram_depth = 8192;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a28.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a28.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a28.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cyclone10lp_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "C:/RISCV/kyogenrv/fpga/kyogenrv_top.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "kyogenrv_fpga_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_63i1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 13;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 8191;
defparam ram_block1a29.port_a_logical_ram_depth = 8192;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a29.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a29.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a29.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

endmodule

module kyogenrv_fpga_kyogenrv_fpga_pio_0 (
	data_out_16,
	data_out_17,
	data_out_18,
	data_out_19,
	data_out_20,
	data_out_21,
	data_out_22,
	data_out_23,
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	data_out_9,
	data_out_10,
	data_out_11,
	data_out_12,
	data_out_13,
	data_out_14,
	data_out_15,
	data_out_24,
	data_out_25,
	data_out_26,
	data_out_27,
	data_out_28,
	data_out_29,
	data_out_30,
	data_out_31,
	mem_alu_out_1,
	mem_alu_out_0,
	wait_latency_counter_0,
	mem_ctrl_mem_wr10,
	wait_latency_counter_1,
	reset_n,
	mem_rs_1_0,
	Equal68,
	Equal73,
	writedata,
	mem_alu_out_2,
	mem_alu_out_3,
	mem_rs_1_1,
	mem_rs_1_2,
	mem_rs_1_3,
	mem_rs_1_4,
	mem_rs_1_5,
	mem_rs_1_6,
	mem_rs_1_7,
	mem_rs_1_8,
	data_out_121,
	mem_rs_1_9,
	mem_rs_1_10,
	mem_rs_1_11,
	mem_rs_1_12,
	mem_rs_1_13,
	mem_rs_1_14,
	mem_rs_1_15,
	mem_rs_1_16,
	data_out_171,
	mem_rs_1_17,
	mem_rs_1_18,
	mem_rs_1_19,
	mem_rs_1_20,
	mem_rs_1_21,
	mem_rs_1_22,
	mem_rs_1_23,
	data_out_271,
	readdata_1,
	readdata_0,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	readdata_8,
	readdata_9,
	readdata_10,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_17,
	readdata_18,
	readdata_19,
	readdata_4,
	readdata_2,
	readdata_3,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_20,
	readdata_21,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_27,
	_GEN_73_0,
	clk)/* synthesis synthesis_greybox=0 */;
output 	data_out_16;
output 	data_out_17;
output 	data_out_18;
output 	data_out_19;
output 	data_out_20;
output 	data_out_21;
output 	data_out_22;
output 	data_out_23;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
output 	data_out_8;
output 	data_out_9;
output 	data_out_10;
output 	data_out_11;
output 	data_out_12;
output 	data_out_13;
output 	data_out_14;
output 	data_out_15;
output 	data_out_24;
output 	data_out_25;
output 	data_out_26;
output 	data_out_27;
output 	data_out_28;
output 	data_out_29;
output 	data_out_30;
output 	data_out_31;
input 	mem_alu_out_1;
input 	mem_alu_out_0;
input 	wait_latency_counter_0;
input 	mem_ctrl_mem_wr10;
input 	wait_latency_counter_1;
input 	reset_n;
input 	mem_rs_1_0;
input 	Equal68;
input 	Equal73;
input 	[31:0] writedata;
input 	mem_alu_out_2;
input 	mem_alu_out_3;
input 	mem_rs_1_1;
input 	mem_rs_1_2;
input 	mem_rs_1_3;
input 	mem_rs_1_4;
input 	mem_rs_1_5;
input 	mem_rs_1_6;
input 	mem_rs_1_7;
input 	mem_rs_1_8;
output 	data_out_121;
input 	mem_rs_1_9;
input 	mem_rs_1_10;
input 	mem_rs_1_11;
input 	mem_rs_1_12;
input 	mem_rs_1_13;
input 	mem_rs_1_14;
input 	mem_rs_1_15;
input 	mem_rs_1_16;
output 	data_out_171;
input 	mem_rs_1_17;
input 	mem_rs_1_18;
input 	mem_rs_1_19;
input 	mem_rs_1_20;
input 	mem_rs_1_21;
input 	mem_rs_1_22;
input 	mem_rs_1_23;
output 	data_out_271;
output 	readdata_1;
output 	readdata_0;
output 	readdata_28;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
output 	readdata_8;
output 	readdata_9;
output 	readdata_10;
output 	readdata_11;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
output 	readdata_15;
output 	readdata_16;
output 	readdata_17;
output 	readdata_18;
output 	readdata_19;
output 	readdata_4;
output 	readdata_2;
output 	readdata_3;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_20;
output 	readdata_21;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_27;
input 	_GEN_73_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_out[17]~10_combout ;
wire \data_out[16]~0_combout ;
wire \data_out[17]~12_combout ;
wire \always0~0_combout ;
wire \always0~1_combout ;
wire \data_out[17]~1_combout ;
wire \data_out[18]~2_combout ;
wire \data_out[19]~3_combout ;
wire \data_out[20]~4_combout ;
wire \data_out[21]~5_combout ;
wire \data_out[22]~6_combout ;
wire \data_out[23]~7_combout ;
wire \data_out[12]~8_combout ;


dffeas \data_out[16] (
	.clk(clk),
	.d(\data_out[16]~0_combout ),
	.asdata(mem_rs_1_16),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\data_out[17]~12_combout ),
	.sload(_GEN_73_0),
	.ena(\always0~1_combout ),
	.q(data_out_16),
	.prn(vcc));
defparam \data_out[16] .is_wysiwyg = "true";
defparam \data_out[16] .power_up = "low";

dffeas \data_out[17] (
	.clk(clk),
	.d(\data_out[17]~1_combout ),
	.asdata(mem_rs_1_17),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\data_out[17]~12_combout ),
	.sload(_GEN_73_0),
	.ena(\always0~1_combout ),
	.q(data_out_17),
	.prn(vcc));
defparam \data_out[17] .is_wysiwyg = "true";
defparam \data_out[17] .power_up = "low";

dffeas \data_out[18] (
	.clk(clk),
	.d(\data_out[18]~2_combout ),
	.asdata(mem_rs_1_18),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\data_out[17]~12_combout ),
	.sload(_GEN_73_0),
	.ena(\always0~1_combout ),
	.q(data_out_18),
	.prn(vcc));
defparam \data_out[18] .is_wysiwyg = "true";
defparam \data_out[18] .power_up = "low";

dffeas \data_out[19] (
	.clk(clk),
	.d(\data_out[19]~3_combout ),
	.asdata(mem_rs_1_19),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\data_out[17]~12_combout ),
	.sload(_GEN_73_0),
	.ena(\always0~1_combout ),
	.q(data_out_19),
	.prn(vcc));
defparam \data_out[19] .is_wysiwyg = "true";
defparam \data_out[19] .power_up = "low";

dffeas \data_out[20] (
	.clk(clk),
	.d(\data_out[20]~4_combout ),
	.asdata(mem_rs_1_20),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\data_out[17]~12_combout ),
	.sload(_GEN_73_0),
	.ena(\always0~1_combout ),
	.q(data_out_20),
	.prn(vcc));
defparam \data_out[20] .is_wysiwyg = "true";
defparam \data_out[20] .power_up = "low";

dffeas \data_out[21] (
	.clk(clk),
	.d(\data_out[21]~5_combout ),
	.asdata(mem_rs_1_21),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\data_out[17]~12_combout ),
	.sload(_GEN_73_0),
	.ena(\always0~1_combout ),
	.q(data_out_21),
	.prn(vcc));
defparam \data_out[21] .is_wysiwyg = "true";
defparam \data_out[21] .power_up = "low";

dffeas \data_out[22] (
	.clk(clk),
	.d(\data_out[22]~6_combout ),
	.asdata(mem_rs_1_22),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\data_out[17]~12_combout ),
	.sload(_GEN_73_0),
	.ena(\always0~1_combout ),
	.q(data_out_22),
	.prn(vcc));
defparam \data_out[22] .is_wysiwyg = "true";
defparam \data_out[22] .power_up = "low";

dffeas \data_out[23] (
	.clk(clk),
	.d(\data_out[23]~7_combout ),
	.asdata(mem_rs_1_23),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\data_out[17]~12_combout ),
	.sload(_GEN_73_0),
	.ena(\always0~1_combout ),
	.q(data_out_23),
	.prn(vcc));
defparam \data_out[23] .is_wysiwyg = "true";
defparam \data_out[23] .power_up = "low";

dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

dffeas \data_out[8] (
	.clk(clk),
	.d(writedata[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_8),
	.prn(vcc));
defparam \data_out[8] .is_wysiwyg = "true";
defparam \data_out[8] .power_up = "low";

dffeas \data_out[9] (
	.clk(clk),
	.d(writedata[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_9),
	.prn(vcc));
defparam \data_out[9] .is_wysiwyg = "true";
defparam \data_out[9] .power_up = "low";

dffeas \data_out[10] (
	.clk(clk),
	.d(writedata[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_10),
	.prn(vcc));
defparam \data_out[10] .is_wysiwyg = "true";
defparam \data_out[10] .power_up = "low";

dffeas \data_out[11] (
	.clk(clk),
	.d(writedata[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_11),
	.prn(vcc));
defparam \data_out[11] .is_wysiwyg = "true";
defparam \data_out[11] .power_up = "low";

dffeas \data_out[12] (
	.clk(clk),
	.d(writedata[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_12),
	.prn(vcc));
defparam \data_out[12] .is_wysiwyg = "true";
defparam \data_out[12] .power_up = "low";

dffeas \data_out[13] (
	.clk(clk),
	.d(writedata[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_13),
	.prn(vcc));
defparam \data_out[13] .is_wysiwyg = "true";
defparam \data_out[13] .power_up = "low";

dffeas \data_out[14] (
	.clk(clk),
	.d(writedata[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_14),
	.prn(vcc));
defparam \data_out[14] .is_wysiwyg = "true";
defparam \data_out[14] .power_up = "low";

dffeas \data_out[15] (
	.clk(clk),
	.d(writedata[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_15),
	.prn(vcc));
defparam \data_out[15] .is_wysiwyg = "true";
defparam \data_out[15] .power_up = "low";

dffeas \data_out[24] (
	.clk(clk),
	.d(writedata[24]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_24),
	.prn(vcc));
defparam \data_out[24] .is_wysiwyg = "true";
defparam \data_out[24] .power_up = "low";

dffeas \data_out[25] (
	.clk(clk),
	.d(writedata[25]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_25),
	.prn(vcc));
defparam \data_out[25] .is_wysiwyg = "true";
defparam \data_out[25] .power_up = "low";

dffeas \data_out[26] (
	.clk(clk),
	.d(writedata[26]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_26),
	.prn(vcc));
defparam \data_out[26] .is_wysiwyg = "true";
defparam \data_out[26] .power_up = "low";

dffeas \data_out[27] (
	.clk(clk),
	.d(writedata[27]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_27),
	.prn(vcc));
defparam \data_out[27] .is_wysiwyg = "true";
defparam \data_out[27] .power_up = "low";

dffeas \data_out[28] (
	.clk(clk),
	.d(writedata[28]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_28),
	.prn(vcc));
defparam \data_out[28] .is_wysiwyg = "true";
defparam \data_out[28] .power_up = "low";

dffeas \data_out[29] (
	.clk(clk),
	.d(writedata[29]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_29),
	.prn(vcc));
defparam \data_out[29] .is_wysiwyg = "true";
defparam \data_out[29] .power_up = "low";

dffeas \data_out[30] (
	.clk(clk),
	.d(writedata[30]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_30),
	.prn(vcc));
defparam \data_out[30] .is_wysiwyg = "true";
defparam \data_out[30] .power_up = "low";

dffeas \data_out[31] (
	.clk(clk),
	.d(writedata[31]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_31),
	.prn(vcc));
defparam \data_out[31] .is_wysiwyg = "true";
defparam \data_out[31] .power_up = "low";

cyclone10lp_lcell_comb \data_out[12]~9 (
	.dataa(\data_out[12]~8_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_ctrl_mem_wr10),
	.cin(gnd),
	.combout(data_out_121),
	.cout());
defparam \data_out[12]~9 .lut_mask = 16'hAAFF;
defparam \data_out[12]~9 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[17]~11 (
	.dataa(mem_alu_out_0),
	.datab(Equal68),
	.datac(Equal73),
	.datad(gnd),
	.cin(gnd),
	.combout(data_out_171),
	.cout());
defparam \data_out[17]~11 .lut_mask = 16'hA8A8;
defparam \data_out[17]~11 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[27]~13 (
	.dataa(mem_alu_out_0),
	.datab(mem_alu_out_1),
	.datac(Equal68),
	.datad(Equal73),
	.cin(gnd),
	.combout(data_out_271),
	.cout());
defparam \data_out[27]~13 .lut_mask = 16'h999F;
defparam \data_out[27]~13 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[1] (
	.dataa(data_out_1),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1] .lut_mask = 16'h000A;
defparam \readdata[1] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[0] (
	.dataa(data_out_0),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0] .lut_mask = 16'h000A;
defparam \readdata[0] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[28] (
	.dataa(data_out_28),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_28),
	.cout());
defparam \readdata[28] .lut_mask = 16'h000A;
defparam \readdata[28] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[29] (
	.dataa(data_out_29),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_29),
	.cout());
defparam \readdata[29] .lut_mask = 16'h000A;
defparam \readdata[29] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[30] (
	.dataa(data_out_30),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_30),
	.cout());
defparam \readdata[30] .lut_mask = 16'h000A;
defparam \readdata[30] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[31] (
	.dataa(data_out_31),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_31),
	.cout());
defparam \readdata[31] .lut_mask = 16'h000A;
defparam \readdata[31] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[8] (
	.dataa(data_out_8),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_8),
	.cout());
defparam \readdata[8] .lut_mask = 16'h000A;
defparam \readdata[8] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[9] (
	.dataa(data_out_9),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_9),
	.cout());
defparam \readdata[9] .lut_mask = 16'h000A;
defparam \readdata[9] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[10] (
	.dataa(data_out_10),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_10),
	.cout());
defparam \readdata[10] .lut_mask = 16'h000A;
defparam \readdata[10] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[11] (
	.dataa(data_out_11),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_11),
	.cout());
defparam \readdata[11] .lut_mask = 16'h000A;
defparam \readdata[11] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[12] (
	.dataa(data_out_12),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_12),
	.cout());
defparam \readdata[12] .lut_mask = 16'h000A;
defparam \readdata[12] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[13] (
	.dataa(data_out_13),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_13),
	.cout());
defparam \readdata[13] .lut_mask = 16'h000A;
defparam \readdata[13] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[14] (
	.dataa(data_out_14),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_14),
	.cout());
defparam \readdata[14] .lut_mask = 16'h000A;
defparam \readdata[14] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[15] (
	.dataa(data_out_15),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_15),
	.cout());
defparam \readdata[15] .lut_mask = 16'h000A;
defparam \readdata[15] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[16] (
	.dataa(data_out_16),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_16),
	.cout());
defparam \readdata[16] .lut_mask = 16'h000A;
defparam \readdata[16] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[17] (
	.dataa(data_out_17),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_17),
	.cout());
defparam \readdata[17] .lut_mask = 16'h000A;
defparam \readdata[17] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[18] (
	.dataa(data_out_18),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_18),
	.cout());
defparam \readdata[18] .lut_mask = 16'h000A;
defparam \readdata[18] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[19] (
	.dataa(data_out_19),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_19),
	.cout());
defparam \readdata[19] .lut_mask = 16'h000A;
defparam \readdata[19] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[4] (
	.dataa(data_out_4),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_4),
	.cout());
defparam \readdata[4] .lut_mask = 16'h000A;
defparam \readdata[4] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[2] (
	.dataa(data_out_2),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_2),
	.cout());
defparam \readdata[2] .lut_mask = 16'h000A;
defparam \readdata[2] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[3] (
	.dataa(data_out_3),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_3),
	.cout());
defparam \readdata[3] .lut_mask = 16'h000A;
defparam \readdata[3] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[5] (
	.dataa(data_out_5),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_5),
	.cout());
defparam \readdata[5] .lut_mask = 16'h000A;
defparam \readdata[5] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[6] (
	.dataa(data_out_6),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_6),
	.cout());
defparam \readdata[6] .lut_mask = 16'h000A;
defparam \readdata[6] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[7] (
	.dataa(data_out_7),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_7),
	.cout());
defparam \readdata[7] .lut_mask = 16'h000A;
defparam \readdata[7] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[20] (
	.dataa(data_out_20),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_20),
	.cout());
defparam \readdata[20] .lut_mask = 16'h000A;
defparam \readdata[20] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[21] (
	.dataa(data_out_21),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_21),
	.cout());
defparam \readdata[21] .lut_mask = 16'h000A;
defparam \readdata[21] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[22] (
	.dataa(data_out_22),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_22),
	.cout());
defparam \readdata[22] .lut_mask = 16'h000A;
defparam \readdata[22] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[23] (
	.dataa(data_out_23),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_23),
	.cout());
defparam \readdata[23] .lut_mask = 16'h000A;
defparam \readdata[23] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[24] (
	.dataa(data_out_24),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_24),
	.cout());
defparam \readdata[24] .lut_mask = 16'h000A;
defparam \readdata[24] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[25] (
	.dataa(data_out_25),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_25),
	.cout());
defparam \readdata[25] .lut_mask = 16'h000A;
defparam \readdata[25] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[26] (
	.dataa(data_out_26),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_26),
	.cout());
defparam \readdata[26] .lut_mask = 16'h000A;
defparam \readdata[26] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \readdata[27] (
	.dataa(data_out_27),
	.datab(gnd),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(readdata_27),
	.cout());
defparam \readdata[27] .lut_mask = 16'h000A;
defparam \readdata[27] .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[17]~10 (
	.dataa(mem_alu_out_1),
	.datab(gnd),
	.datac(mem_alu_out_0),
	.datad(Equal68),
	.cin(gnd),
	.combout(\data_out[17]~10_combout ),
	.cout());
defparam \data_out[17]~10 .lut_mask = 16'hAFFF;
defparam \data_out[17]~10 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[16]~0 (
	.dataa(mem_rs_1_8),
	.datab(mem_rs_1_0),
	.datac(gnd),
	.datad(\data_out[17]~10_combout ),
	.cin(gnd),
	.combout(\data_out[16]~0_combout ),
	.cout());
defparam \data_out[16]~0 .lut_mask = 16'hCCAA;
defparam \data_out[16]~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[17]~12 (
	.dataa(\data_out[17]~10_combout ),
	.datab(data_out_171),
	.datac(gnd),
	.datad(mem_ctrl_mem_wr10),
	.cin(gnd),
	.combout(\data_out[17]~12_combout ),
	.cout());
defparam \data_out[17]~12 .lut_mask = 16'h88FF;
defparam \data_out[17]~12 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \always0~0 (
	.dataa(wait_latency_counter_0),
	.datab(wait_latency_counter_1),
	.datac(mem_alu_out_2),
	.datad(mem_alu_out_3),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'h0001;
defparam \always0~0 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \always0~1 (
	.dataa(mem_ctrl_mem_wr10),
	.datab(\always0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
defparam \always0~1 .lut_mask = 16'h8888;
defparam \always0~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[17]~1 (
	.dataa(mem_rs_1_9),
	.datab(mem_rs_1_1),
	.datac(gnd),
	.datad(\data_out[17]~10_combout ),
	.cin(gnd),
	.combout(\data_out[17]~1_combout ),
	.cout());
defparam \data_out[17]~1 .lut_mask = 16'hCCAA;
defparam \data_out[17]~1 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[18]~2 (
	.dataa(mem_rs_1_10),
	.datab(mem_rs_1_2),
	.datac(gnd),
	.datad(\data_out[17]~10_combout ),
	.cin(gnd),
	.combout(\data_out[18]~2_combout ),
	.cout());
defparam \data_out[18]~2 .lut_mask = 16'hCCAA;
defparam \data_out[18]~2 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[19]~3 (
	.dataa(mem_rs_1_11),
	.datab(mem_rs_1_3),
	.datac(gnd),
	.datad(\data_out[17]~10_combout ),
	.cin(gnd),
	.combout(\data_out[19]~3_combout ),
	.cout());
defparam \data_out[19]~3 .lut_mask = 16'hCCAA;
defparam \data_out[19]~3 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[20]~4 (
	.dataa(mem_rs_1_12),
	.datab(mem_rs_1_4),
	.datac(gnd),
	.datad(\data_out[17]~10_combout ),
	.cin(gnd),
	.combout(\data_out[20]~4_combout ),
	.cout());
defparam \data_out[20]~4 .lut_mask = 16'hCCAA;
defparam \data_out[20]~4 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[21]~5 (
	.dataa(mem_rs_1_13),
	.datab(mem_rs_1_5),
	.datac(gnd),
	.datad(\data_out[17]~10_combout ),
	.cin(gnd),
	.combout(\data_out[21]~5_combout ),
	.cout());
defparam \data_out[21]~5 .lut_mask = 16'hCCAA;
defparam \data_out[21]~5 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[22]~6 (
	.dataa(mem_rs_1_14),
	.datab(mem_rs_1_6),
	.datac(gnd),
	.datad(\data_out[17]~10_combout ),
	.cin(gnd),
	.combout(\data_out[22]~6_combout ),
	.cout());
defparam \data_out[22]~6 .lut_mask = 16'hCCAA;
defparam \data_out[22]~6 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[23]~7 (
	.dataa(mem_rs_1_15),
	.datab(mem_rs_1_7),
	.datac(gnd),
	.datad(\data_out[17]~10_combout ),
	.cin(gnd),
	.combout(\data_out[23]~7_combout ),
	.cout());
defparam \data_out[23]~7 .lut_mask = 16'hCCAA;
defparam \data_out[23]~7 .sum_lutc_input = "datac";

cyclone10lp_lcell_comb \data_out[12]~8 (
	.dataa(mem_alu_out_1),
	.datab(Equal73),
	.datac(mem_alu_out_0),
	.datad(Equal68),
	.cin(gnd),
	.combout(\data_out[12]~8_combout ),
	.cout());
defparam \data_out[12]~8 .lut_mask = 16'hAAC8;
defparam \data_out[12]~8 .sum_lutc_input = "datac";

endmodule
