// kyogenrv_fpga.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module kyogenrv_fpga (
		input  wire        clk_clk,                          //                       clk.clk
		output wire [31:0] kyogenrv_0_counter_readdata,      //        kyogenrv_0_counter.readdata
		output wire [31:0] pio_0_external_connection_export, // pio_0_external_connection.export
		input  wire        reset_reset_n                     //                     reset.reset_n
	);

	wire  [31:0] kyogenrv_0_avalon_data_master_readdata;             // mm_interconnect_0:KyogenRV_0_avalon_data_master_readdata -> KyogenRV_0:r_dmem_data
	wire         kyogenrv_0_avalon_data_master_waitrequest;          // mm_interconnect_0:KyogenRV_0_avalon_data_master_waitrequest -> KyogenRV_0:dmem_waitrequest
	wire   [3:0] kyogenrv_0_avalon_data_master_byteenable;           // KyogenRV_0:w_dmem_data_byteenable -> mm_interconnect_0:KyogenRV_0_avalon_data_master_byteenable
	wire  [31:0] kyogenrv_0_avalon_data_master_address;              // KyogenRV_0:dmem_addr -> mm_interconnect_0:KyogenRV_0_avalon_data_master_address
	wire         kyogenrv_0_avalon_data_master_read;                 // KyogenRV_0:r_dmem_data_req -> mm_interconnect_0:KyogenRV_0_avalon_data_master_read
	wire         kyogenrv_0_avalon_data_master_readdatavalid;        // mm_interconnect_0:KyogenRV_0_avalon_data_master_readdatavalid -> KyogenRV_0:r_dmem_data_ack
	wire  [31:0] kyogenrv_0_avalon_data_master_writedata;            // KyogenRV_0:w_dmem_data -> mm_interconnect_0:KyogenRV_0_avalon_data_master_writedata
	wire         kyogenrv_0_avalon_data_master_write;                // KyogenRV_0:w_dmem_data_req -> mm_interconnect_0:KyogenRV_0_avalon_data_master_write
	wire         mm_interconnect_0_pio_0_s1_chipselect;              // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                 // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;                   // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;               // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire  [31:0] kyogenrv_0_avalon_instruction_master_readdata;      // mm_interconnect_1:KyogenRV_0_avalon_instruction_master_readdata -> KyogenRV_0:r_imem_data
	wire         kyogenrv_0_avalon_instruction_master_waitrequest;   // mm_interconnect_1:KyogenRV_0_avalon_instruction_master_waitrequest -> KyogenRV_0:imem_waitrequest
	wire   [3:0] kyogenrv_0_avalon_instruction_master_byteenable;    // KyogenRV_0:w_imem_data_byteenable -> mm_interconnect_1:KyogenRV_0_avalon_instruction_master_byteenable
	wire  [31:0] kyogenrv_0_avalon_instruction_master_address;       // KyogenRV_0:imem_addr -> mm_interconnect_1:KyogenRV_0_avalon_instruction_master_address
	wire         kyogenrv_0_avalon_instruction_master_read;          // KyogenRV_0:r_imem_data_req -> mm_interconnect_1:KyogenRV_0_avalon_instruction_master_read
	wire         kyogenrv_0_avalon_instruction_master_readdatavalid; // mm_interconnect_1:KyogenRV_0_avalon_instruction_master_readdatavalid -> KyogenRV_0:r_imem_data_ack
	wire  [31:0] kyogenrv_0_avalon_instruction_master_writedata;     // KyogenRV_0:w_imem_data -> mm_interconnect_1:KyogenRV_0_avalon_instruction_master_writedata
	wire         kyogenrv_0_avalon_instruction_master_write;         // KyogenRV_0:w_imem_data_req -> mm_interconnect_1:KyogenRV_0_avalon_instruction_master_write
	wire         mm_interconnect_1_onchip_memory2_0_s1_chipselect;   // mm_interconnect_1:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s1_readdata;     // onchip_memory2_0:readdata -> mm_interconnect_1:onchip_memory2_0_s1_readdata
	wire  [12:0] mm_interconnect_1_onchip_memory2_0_s1_address;      // mm_interconnect_1:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_1_onchip_memory2_0_s1_byteenable;   // mm_interconnect_1:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_1_onchip_memory2_0_s1_write;        // mm_interconnect_1:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s1_writedata;    // mm_interconnect_1:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_1_onchip_memory2_0_s1_clken;        // mm_interconnect_1:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         rst_controller_reset_out_reset;                     // rst_controller:reset_out -> [KyogenRV_0:reset, mm_interconnect_0:KyogenRV_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:KyogenRV_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, pio_0:reset_n]

	kyogenrv_fpga_KyogenRV_0 kyogenrv_0 (
		.reset                  (rst_controller_reset_out_reset),                     //                     reset.reset
		.clock                  (clk_clk),                                            //                clock_sink.clk
		.r_imem_data_ack        (kyogenrv_0_avalon_instruction_master_readdatavalid), // avalon_instruction_master.readdatavalid
		.r_imem_data            (kyogenrv_0_avalon_instruction_master_readdata),      //                          .readdata
		.w_imem_data            (kyogenrv_0_avalon_instruction_master_writedata),     //                          .writedata
		.w_imem_data_byteenable (kyogenrv_0_avalon_instruction_master_byteenable),    //                          .byteenable
		.imem_addr              (kyogenrv_0_avalon_instruction_master_address),       //                          .address
		.imem_waitrequest       (kyogenrv_0_avalon_instruction_master_waitrequest),   //                          .waitrequest
		.r_imem_data_req        (kyogenrv_0_avalon_instruction_master_read),          //                          .read
		.w_imem_data_req        (kyogenrv_0_avalon_instruction_master_write),         //                          .write
		.w_dmem_data            (kyogenrv_0_avalon_data_master_writedata),            //        avalon_data_master.writedata
		.w_dmem_data_byteenable (kyogenrv_0_avalon_data_master_byteenable),           //                          .byteenable
		.r_dmem_data_ack        (kyogenrv_0_avalon_data_master_readdatavalid),        //                          .readdatavalid
		.dmem_addr              (kyogenrv_0_avalon_data_master_address),              //                          .address
		.r_dmem_data            (kyogenrv_0_avalon_data_master_readdata),             //                          .readdata
		.dmem_waitrequest       (kyogenrv_0_avalon_data_master_waitrequest),          //                          .waitrequest
		.r_dmem_data_req        (kyogenrv_0_avalon_data_master_read),                 //                          .read
		.w_dmem_data_req        (kyogenrv_0_avalon_data_master_write),                //                          .write
		.pc_counter             (kyogenrv_0_counter_readdata)                         //                   counter.readdata
	);

	kyogenrv_fpga_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_1_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_1_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (1'b0),                                             // (terminated)
		.freeze     (1'b0)                                              // (terminated)
	);

	kyogenrv_fpga_pio_0 pio_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (pio_0_external_connection_export)       // external_connection.export
	);

	kyogenrv_fpga_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                (clk_clk),                                     //                              clk_0_clk.clk
		.KyogenRV_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),              // KyogenRV_0_reset_reset_bridge_in_reset.reset
		.KyogenRV_0_avalon_data_master_address        (kyogenrv_0_avalon_data_master_address),       //          KyogenRV_0_avalon_data_master.address
		.KyogenRV_0_avalon_data_master_waitrequest    (kyogenrv_0_avalon_data_master_waitrequest),   //                                       .waitrequest
		.KyogenRV_0_avalon_data_master_byteenable     (kyogenrv_0_avalon_data_master_byteenable),    //                                       .byteenable
		.KyogenRV_0_avalon_data_master_read           (kyogenrv_0_avalon_data_master_read),          //                                       .read
		.KyogenRV_0_avalon_data_master_readdata       (kyogenrv_0_avalon_data_master_readdata),      //                                       .readdata
		.KyogenRV_0_avalon_data_master_readdatavalid  (kyogenrv_0_avalon_data_master_readdatavalid), //                                       .readdatavalid
		.KyogenRV_0_avalon_data_master_write          (kyogenrv_0_avalon_data_master_write),         //                                       .write
		.KyogenRV_0_avalon_data_master_writedata      (kyogenrv_0_avalon_data_master_writedata),     //                                       .writedata
		.pio_0_s1_address                             (mm_interconnect_0_pio_0_s1_address),          //                               pio_0_s1.address
		.pio_0_s1_write                               (mm_interconnect_0_pio_0_s1_write),            //                                       .write
		.pio_0_s1_readdata                            (mm_interconnect_0_pio_0_s1_readdata),         //                                       .readdata
		.pio_0_s1_writedata                           (mm_interconnect_0_pio_0_s1_writedata),        //                                       .writedata
		.pio_0_s1_chipselect                          (mm_interconnect_0_pio_0_s1_chipselect)        //                                       .chipselect
	);

	kyogenrv_fpga_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                      (clk_clk),                                            //                              clk_0_clk.clk
		.KyogenRV_0_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                     // KyogenRV_0_reset_reset_bridge_in_reset.reset
		.KyogenRV_0_avalon_instruction_master_address       (kyogenrv_0_avalon_instruction_master_address),       //   KyogenRV_0_avalon_instruction_master.address
		.KyogenRV_0_avalon_instruction_master_waitrequest   (kyogenrv_0_avalon_instruction_master_waitrequest),   //                                       .waitrequest
		.KyogenRV_0_avalon_instruction_master_byteenable    (kyogenrv_0_avalon_instruction_master_byteenable),    //                                       .byteenable
		.KyogenRV_0_avalon_instruction_master_read          (kyogenrv_0_avalon_instruction_master_read),          //                                       .read
		.KyogenRV_0_avalon_instruction_master_readdata      (kyogenrv_0_avalon_instruction_master_readdata),      //                                       .readdata
		.KyogenRV_0_avalon_instruction_master_readdatavalid (kyogenrv_0_avalon_instruction_master_readdatavalid), //                                       .readdatavalid
		.KyogenRV_0_avalon_instruction_master_write         (kyogenrv_0_avalon_instruction_master_write),         //                                       .write
		.KyogenRV_0_avalon_instruction_master_writedata     (kyogenrv_0_avalon_instruction_master_writedata),     //                                       .writedata
		.onchip_memory2_0_s1_address                        (mm_interconnect_1_onchip_memory2_0_s1_address),      //                    onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                          (mm_interconnect_1_onchip_memory2_0_s1_write),        //                                       .write
		.onchip_memory2_0_s1_readdata                       (mm_interconnect_1_onchip_memory2_0_s1_readdata),     //                                       .readdata
		.onchip_memory2_0_s1_writedata                      (mm_interconnect_1_onchip_memory2_0_s1_writedata),    //                                       .writedata
		.onchip_memory2_0_s1_byteenable                     (mm_interconnect_1_onchip_memory2_0_s1_byteenable),   //                                       .byteenable
		.onchip_memory2_0_s1_chipselect                     (mm_interconnect_1_onchip_memory2_0_s1_chipselect),   //                                       .chipselect
		.onchip_memory2_0_s1_clken                          (mm_interconnect_1_onchip_memory2_0_s1_clken)         //                                       .clken
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
